
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
-- All structs defined in C code

package c_structs_pkg is
subtype uint1_t is unsigned(0 downto 0);
constant uint1_t_SLV_LEN : integer := 1;
function uint1_t_to_slv(x : uint1_t) return std_logic_vector;
function slv_to_uint1_t(x : std_logic_vector) return uint1_t;
subtype uint2_t is unsigned(1 downto 0);
constant uint2_t_SLV_LEN : integer := 2;
function uint2_t_to_slv(x : uint2_t) return std_logic_vector;
function slv_to_uint2_t(x : std_logic_vector) return uint2_t;
subtype int2_t is signed(1 downto 0);
constant int2_t_SLV_LEN : integer := 2;
function int2_t_to_slv(x : int2_t) return std_logic_vector;
function slv_to_int2_t(x : std_logic_vector) return int2_t;
subtype uint3_t is unsigned(2 downto 0);
constant uint3_t_SLV_LEN : integer := 3;
function uint3_t_to_slv(x : uint3_t) return std_logic_vector;
function slv_to_uint3_t(x : std_logic_vector) return uint3_t;
subtype int3_t is signed(2 downto 0);
constant int3_t_SLV_LEN : integer := 3;
function int3_t_to_slv(x : int3_t) return std_logic_vector;
function slv_to_int3_t(x : std_logic_vector) return int3_t;
subtype uint4_t is unsigned(3 downto 0);
constant uint4_t_SLV_LEN : integer := 4;
function uint4_t_to_slv(x : uint4_t) return std_logic_vector;
function slv_to_uint4_t(x : std_logic_vector) return uint4_t;
subtype int4_t is signed(3 downto 0);
constant int4_t_SLV_LEN : integer := 4;
function int4_t_to_slv(x : int4_t) return std_logic_vector;
function slv_to_int4_t(x : std_logic_vector) return int4_t;
subtype uint5_t is unsigned(4 downto 0);
constant uint5_t_SLV_LEN : integer := 5;
function uint5_t_to_slv(x : uint5_t) return std_logic_vector;
function slv_to_uint5_t(x : std_logic_vector) return uint5_t;
subtype int5_t is signed(4 downto 0);
constant int5_t_SLV_LEN : integer := 5;
function int5_t_to_slv(x : int5_t) return std_logic_vector;
function slv_to_int5_t(x : std_logic_vector) return int5_t;
subtype uint6_t is unsigned(5 downto 0);
constant uint6_t_SLV_LEN : integer := 6;
function uint6_t_to_slv(x : uint6_t) return std_logic_vector;
function slv_to_uint6_t(x : std_logic_vector) return uint6_t;
subtype int6_t is signed(5 downto 0);
constant int6_t_SLV_LEN : integer := 6;
function int6_t_to_slv(x : int6_t) return std_logic_vector;
function slv_to_int6_t(x : std_logic_vector) return int6_t;
subtype uint7_t is unsigned(6 downto 0);
constant uint7_t_SLV_LEN : integer := 7;
function uint7_t_to_slv(x : uint7_t) return std_logic_vector;
function slv_to_uint7_t(x : std_logic_vector) return uint7_t;
subtype int7_t is signed(6 downto 0);
constant int7_t_SLV_LEN : integer := 7;
function int7_t_to_slv(x : int7_t) return std_logic_vector;
function slv_to_int7_t(x : std_logic_vector) return int7_t;
subtype uint8_t is unsigned(7 downto 0);
constant uint8_t_SLV_LEN : integer := 8;
function uint8_t_to_slv(x : uint8_t) return std_logic_vector;
function slv_to_uint8_t(x : std_logic_vector) return uint8_t;
subtype int8_t is signed(7 downto 0);
constant int8_t_SLV_LEN : integer := 8;
function int8_t_to_slv(x : int8_t) return std_logic_vector;
function slv_to_int8_t(x : std_logic_vector) return int8_t;
subtype uint9_t is unsigned(8 downto 0);
constant uint9_t_SLV_LEN : integer := 9;
function uint9_t_to_slv(x : uint9_t) return std_logic_vector;
function slv_to_uint9_t(x : std_logic_vector) return uint9_t;
subtype int9_t is signed(8 downto 0);
constant int9_t_SLV_LEN : integer := 9;
function int9_t_to_slv(x : int9_t) return std_logic_vector;
function slv_to_int9_t(x : std_logic_vector) return int9_t;
subtype uint10_t is unsigned(9 downto 0);
constant uint10_t_SLV_LEN : integer := 10;
function uint10_t_to_slv(x : uint10_t) return std_logic_vector;
function slv_to_uint10_t(x : std_logic_vector) return uint10_t;
subtype int10_t is signed(9 downto 0);
constant int10_t_SLV_LEN : integer := 10;
function int10_t_to_slv(x : int10_t) return std_logic_vector;
function slv_to_int10_t(x : std_logic_vector) return int10_t;
subtype uint11_t is unsigned(10 downto 0);
constant uint11_t_SLV_LEN : integer := 11;
function uint11_t_to_slv(x : uint11_t) return std_logic_vector;
function slv_to_uint11_t(x : std_logic_vector) return uint11_t;
subtype int11_t is signed(10 downto 0);
constant int11_t_SLV_LEN : integer := 11;
function int11_t_to_slv(x : int11_t) return std_logic_vector;
function slv_to_int11_t(x : std_logic_vector) return int11_t;
subtype uint12_t is unsigned(11 downto 0);
constant uint12_t_SLV_LEN : integer := 12;
function uint12_t_to_slv(x : uint12_t) return std_logic_vector;
function slv_to_uint12_t(x : std_logic_vector) return uint12_t;
subtype int12_t is signed(11 downto 0);
constant int12_t_SLV_LEN : integer := 12;
function int12_t_to_slv(x : int12_t) return std_logic_vector;
function slv_to_int12_t(x : std_logic_vector) return int12_t;
subtype uint13_t is unsigned(12 downto 0);
constant uint13_t_SLV_LEN : integer := 13;
function uint13_t_to_slv(x : uint13_t) return std_logic_vector;
function slv_to_uint13_t(x : std_logic_vector) return uint13_t;
subtype int13_t is signed(12 downto 0);
constant int13_t_SLV_LEN : integer := 13;
function int13_t_to_slv(x : int13_t) return std_logic_vector;
function slv_to_int13_t(x : std_logic_vector) return int13_t;
subtype uint14_t is unsigned(13 downto 0);
constant uint14_t_SLV_LEN : integer := 14;
function uint14_t_to_slv(x : uint14_t) return std_logic_vector;
function slv_to_uint14_t(x : std_logic_vector) return uint14_t;
subtype int14_t is signed(13 downto 0);
constant int14_t_SLV_LEN : integer := 14;
function int14_t_to_slv(x : int14_t) return std_logic_vector;
function slv_to_int14_t(x : std_logic_vector) return int14_t;
subtype uint15_t is unsigned(14 downto 0);
constant uint15_t_SLV_LEN : integer := 15;
function uint15_t_to_slv(x : uint15_t) return std_logic_vector;
function slv_to_uint15_t(x : std_logic_vector) return uint15_t;
subtype int15_t is signed(14 downto 0);
constant int15_t_SLV_LEN : integer := 15;
function int15_t_to_slv(x : int15_t) return std_logic_vector;
function slv_to_int15_t(x : std_logic_vector) return int15_t;
subtype uint16_t is unsigned(15 downto 0);
constant uint16_t_SLV_LEN : integer := 16;
function uint16_t_to_slv(x : uint16_t) return std_logic_vector;
function slv_to_uint16_t(x : std_logic_vector) return uint16_t;
subtype int16_t is signed(15 downto 0);
constant int16_t_SLV_LEN : integer := 16;
function int16_t_to_slv(x : int16_t) return std_logic_vector;
function slv_to_int16_t(x : std_logic_vector) return int16_t;
subtype uint17_t is unsigned(16 downto 0);
constant uint17_t_SLV_LEN : integer := 17;
function uint17_t_to_slv(x : uint17_t) return std_logic_vector;
function slv_to_uint17_t(x : std_logic_vector) return uint17_t;
subtype int17_t is signed(16 downto 0);
constant int17_t_SLV_LEN : integer := 17;
function int17_t_to_slv(x : int17_t) return std_logic_vector;
function slv_to_int17_t(x : std_logic_vector) return int17_t;
subtype uint18_t is unsigned(17 downto 0);
constant uint18_t_SLV_LEN : integer := 18;
function uint18_t_to_slv(x : uint18_t) return std_logic_vector;
function slv_to_uint18_t(x : std_logic_vector) return uint18_t;
subtype int18_t is signed(17 downto 0);
constant int18_t_SLV_LEN : integer := 18;
function int18_t_to_slv(x : int18_t) return std_logic_vector;
function slv_to_int18_t(x : std_logic_vector) return int18_t;
subtype uint19_t is unsigned(18 downto 0);
constant uint19_t_SLV_LEN : integer := 19;
function uint19_t_to_slv(x : uint19_t) return std_logic_vector;
function slv_to_uint19_t(x : std_logic_vector) return uint19_t;
subtype int19_t is signed(18 downto 0);
constant int19_t_SLV_LEN : integer := 19;
function int19_t_to_slv(x : int19_t) return std_logic_vector;
function slv_to_int19_t(x : std_logic_vector) return int19_t;
subtype uint20_t is unsigned(19 downto 0);
constant uint20_t_SLV_LEN : integer := 20;
function uint20_t_to_slv(x : uint20_t) return std_logic_vector;
function slv_to_uint20_t(x : std_logic_vector) return uint20_t;
subtype int20_t is signed(19 downto 0);
constant int20_t_SLV_LEN : integer := 20;
function int20_t_to_slv(x : int20_t) return std_logic_vector;
function slv_to_int20_t(x : std_logic_vector) return int20_t;
subtype uint21_t is unsigned(20 downto 0);
constant uint21_t_SLV_LEN : integer := 21;
function uint21_t_to_slv(x : uint21_t) return std_logic_vector;
function slv_to_uint21_t(x : std_logic_vector) return uint21_t;
subtype int21_t is signed(20 downto 0);
constant int21_t_SLV_LEN : integer := 21;
function int21_t_to_slv(x : int21_t) return std_logic_vector;
function slv_to_int21_t(x : std_logic_vector) return int21_t;
subtype uint22_t is unsigned(21 downto 0);
constant uint22_t_SLV_LEN : integer := 22;
function uint22_t_to_slv(x : uint22_t) return std_logic_vector;
function slv_to_uint22_t(x : std_logic_vector) return uint22_t;
subtype int22_t is signed(21 downto 0);
constant int22_t_SLV_LEN : integer := 22;
function int22_t_to_slv(x : int22_t) return std_logic_vector;
function slv_to_int22_t(x : std_logic_vector) return int22_t;
subtype uint23_t is unsigned(22 downto 0);
constant uint23_t_SLV_LEN : integer := 23;
function uint23_t_to_slv(x : uint23_t) return std_logic_vector;
function slv_to_uint23_t(x : std_logic_vector) return uint23_t;
subtype int23_t is signed(22 downto 0);
constant int23_t_SLV_LEN : integer := 23;
function int23_t_to_slv(x : int23_t) return std_logic_vector;
function slv_to_int23_t(x : std_logic_vector) return int23_t;
subtype uint24_t is unsigned(23 downto 0);
constant uint24_t_SLV_LEN : integer := 24;
function uint24_t_to_slv(x : uint24_t) return std_logic_vector;
function slv_to_uint24_t(x : std_logic_vector) return uint24_t;
subtype int24_t is signed(23 downto 0);
constant int24_t_SLV_LEN : integer := 24;
function int24_t_to_slv(x : int24_t) return std_logic_vector;
function slv_to_int24_t(x : std_logic_vector) return int24_t;
subtype uint25_t is unsigned(24 downto 0);
constant uint25_t_SLV_LEN : integer := 25;
function uint25_t_to_slv(x : uint25_t) return std_logic_vector;
function slv_to_uint25_t(x : std_logic_vector) return uint25_t;
subtype int25_t is signed(24 downto 0);
constant int25_t_SLV_LEN : integer := 25;
function int25_t_to_slv(x : int25_t) return std_logic_vector;
function slv_to_int25_t(x : std_logic_vector) return int25_t;
subtype uint26_t is unsigned(25 downto 0);
constant uint26_t_SLV_LEN : integer := 26;
function uint26_t_to_slv(x : uint26_t) return std_logic_vector;
function slv_to_uint26_t(x : std_logic_vector) return uint26_t;
subtype int26_t is signed(25 downto 0);
constant int26_t_SLV_LEN : integer := 26;
function int26_t_to_slv(x : int26_t) return std_logic_vector;
function slv_to_int26_t(x : std_logic_vector) return int26_t;
subtype uint27_t is unsigned(26 downto 0);
constant uint27_t_SLV_LEN : integer := 27;
function uint27_t_to_slv(x : uint27_t) return std_logic_vector;
function slv_to_uint27_t(x : std_logic_vector) return uint27_t;
subtype int27_t is signed(26 downto 0);
constant int27_t_SLV_LEN : integer := 27;
function int27_t_to_slv(x : int27_t) return std_logic_vector;
function slv_to_int27_t(x : std_logic_vector) return int27_t;
subtype uint28_t is unsigned(27 downto 0);
constant uint28_t_SLV_LEN : integer := 28;
function uint28_t_to_slv(x : uint28_t) return std_logic_vector;
function slv_to_uint28_t(x : std_logic_vector) return uint28_t;
subtype int28_t is signed(27 downto 0);
constant int28_t_SLV_LEN : integer := 28;
function int28_t_to_slv(x : int28_t) return std_logic_vector;
function slv_to_int28_t(x : std_logic_vector) return int28_t;
subtype uint29_t is unsigned(28 downto 0);
constant uint29_t_SLV_LEN : integer := 29;
function uint29_t_to_slv(x : uint29_t) return std_logic_vector;
function slv_to_uint29_t(x : std_logic_vector) return uint29_t;
subtype int29_t is signed(28 downto 0);
constant int29_t_SLV_LEN : integer := 29;
function int29_t_to_slv(x : int29_t) return std_logic_vector;
function slv_to_int29_t(x : std_logic_vector) return int29_t;
subtype uint30_t is unsigned(29 downto 0);
constant uint30_t_SLV_LEN : integer := 30;
function uint30_t_to_slv(x : uint30_t) return std_logic_vector;
function slv_to_uint30_t(x : std_logic_vector) return uint30_t;
subtype int30_t is signed(29 downto 0);
constant int30_t_SLV_LEN : integer := 30;
function int30_t_to_slv(x : int30_t) return std_logic_vector;
function slv_to_int30_t(x : std_logic_vector) return int30_t;
subtype uint31_t is unsigned(30 downto 0);
constant uint31_t_SLV_LEN : integer := 31;
function uint31_t_to_slv(x : uint31_t) return std_logic_vector;
function slv_to_uint31_t(x : std_logic_vector) return uint31_t;
subtype int31_t is signed(30 downto 0);
constant int31_t_SLV_LEN : integer := 31;
function int31_t_to_slv(x : int31_t) return std_logic_vector;
function slv_to_int31_t(x : std_logic_vector) return int31_t;
subtype uint32_t is unsigned(31 downto 0);
constant uint32_t_SLV_LEN : integer := 32;
function uint32_t_to_slv(x : uint32_t) return std_logic_vector;
function slv_to_uint32_t(x : std_logic_vector) return uint32_t;
subtype int32_t is signed(31 downto 0);
constant int32_t_SLV_LEN : integer := 32;
function int32_t_to_slv(x : int32_t) return std_logic_vector;
function slv_to_int32_t(x : std_logic_vector) return int32_t;
subtype uint33_t is unsigned(32 downto 0);
constant uint33_t_SLV_LEN : integer := 33;
function uint33_t_to_slv(x : uint33_t) return std_logic_vector;
function slv_to_uint33_t(x : std_logic_vector) return uint33_t;
subtype int33_t is signed(32 downto 0);
constant int33_t_SLV_LEN : integer := 33;
function int33_t_to_slv(x : int33_t) return std_logic_vector;
function slv_to_int33_t(x : std_logic_vector) return int33_t;
subtype uint34_t is unsigned(33 downto 0);
constant uint34_t_SLV_LEN : integer := 34;
function uint34_t_to_slv(x : uint34_t) return std_logic_vector;
function slv_to_uint34_t(x : std_logic_vector) return uint34_t;
subtype int34_t is signed(33 downto 0);
constant int34_t_SLV_LEN : integer := 34;
function int34_t_to_slv(x : int34_t) return std_logic_vector;
function slv_to_int34_t(x : std_logic_vector) return int34_t;
subtype uint35_t is unsigned(34 downto 0);
constant uint35_t_SLV_LEN : integer := 35;
function uint35_t_to_slv(x : uint35_t) return std_logic_vector;
function slv_to_uint35_t(x : std_logic_vector) return uint35_t;
subtype int35_t is signed(34 downto 0);
constant int35_t_SLV_LEN : integer := 35;
function int35_t_to_slv(x : int35_t) return std_logic_vector;
function slv_to_int35_t(x : std_logic_vector) return int35_t;
subtype uint36_t is unsigned(35 downto 0);
constant uint36_t_SLV_LEN : integer := 36;
function uint36_t_to_slv(x : uint36_t) return std_logic_vector;
function slv_to_uint36_t(x : std_logic_vector) return uint36_t;
subtype int36_t is signed(35 downto 0);
constant int36_t_SLV_LEN : integer := 36;
function int36_t_to_slv(x : int36_t) return std_logic_vector;
function slv_to_int36_t(x : std_logic_vector) return int36_t;
subtype uint37_t is unsigned(36 downto 0);
constant uint37_t_SLV_LEN : integer := 37;
function uint37_t_to_slv(x : uint37_t) return std_logic_vector;
function slv_to_uint37_t(x : std_logic_vector) return uint37_t;
subtype int37_t is signed(36 downto 0);
constant int37_t_SLV_LEN : integer := 37;
function int37_t_to_slv(x : int37_t) return std_logic_vector;
function slv_to_int37_t(x : std_logic_vector) return int37_t;
subtype uint38_t is unsigned(37 downto 0);
constant uint38_t_SLV_LEN : integer := 38;
function uint38_t_to_slv(x : uint38_t) return std_logic_vector;
function slv_to_uint38_t(x : std_logic_vector) return uint38_t;
subtype int38_t is signed(37 downto 0);
constant int38_t_SLV_LEN : integer := 38;
function int38_t_to_slv(x : int38_t) return std_logic_vector;
function slv_to_int38_t(x : std_logic_vector) return int38_t;
subtype uint39_t is unsigned(38 downto 0);
constant uint39_t_SLV_LEN : integer := 39;
function uint39_t_to_slv(x : uint39_t) return std_logic_vector;
function slv_to_uint39_t(x : std_logic_vector) return uint39_t;
subtype int39_t is signed(38 downto 0);
constant int39_t_SLV_LEN : integer := 39;
function int39_t_to_slv(x : int39_t) return std_logic_vector;
function slv_to_int39_t(x : std_logic_vector) return int39_t;
subtype uint40_t is unsigned(39 downto 0);
constant uint40_t_SLV_LEN : integer := 40;
function uint40_t_to_slv(x : uint40_t) return std_logic_vector;
function slv_to_uint40_t(x : std_logic_vector) return uint40_t;
subtype int40_t is signed(39 downto 0);
constant int40_t_SLV_LEN : integer := 40;
function int40_t_to_slv(x : int40_t) return std_logic_vector;
function slv_to_int40_t(x : std_logic_vector) return int40_t;
subtype uint41_t is unsigned(40 downto 0);
constant uint41_t_SLV_LEN : integer := 41;
function uint41_t_to_slv(x : uint41_t) return std_logic_vector;
function slv_to_uint41_t(x : std_logic_vector) return uint41_t;
subtype int41_t is signed(40 downto 0);
constant int41_t_SLV_LEN : integer := 41;
function int41_t_to_slv(x : int41_t) return std_logic_vector;
function slv_to_int41_t(x : std_logic_vector) return int41_t;
subtype uint42_t is unsigned(41 downto 0);
constant uint42_t_SLV_LEN : integer := 42;
function uint42_t_to_slv(x : uint42_t) return std_logic_vector;
function slv_to_uint42_t(x : std_logic_vector) return uint42_t;
subtype int42_t is signed(41 downto 0);
constant int42_t_SLV_LEN : integer := 42;
function int42_t_to_slv(x : int42_t) return std_logic_vector;
function slv_to_int42_t(x : std_logic_vector) return int42_t;
subtype uint43_t is unsigned(42 downto 0);
constant uint43_t_SLV_LEN : integer := 43;
function uint43_t_to_slv(x : uint43_t) return std_logic_vector;
function slv_to_uint43_t(x : std_logic_vector) return uint43_t;
subtype int43_t is signed(42 downto 0);
constant int43_t_SLV_LEN : integer := 43;
function int43_t_to_slv(x : int43_t) return std_logic_vector;
function slv_to_int43_t(x : std_logic_vector) return int43_t;
subtype uint44_t is unsigned(43 downto 0);
constant uint44_t_SLV_LEN : integer := 44;
function uint44_t_to_slv(x : uint44_t) return std_logic_vector;
function slv_to_uint44_t(x : std_logic_vector) return uint44_t;
subtype int44_t is signed(43 downto 0);
constant int44_t_SLV_LEN : integer := 44;
function int44_t_to_slv(x : int44_t) return std_logic_vector;
function slv_to_int44_t(x : std_logic_vector) return int44_t;
subtype uint45_t is unsigned(44 downto 0);
constant uint45_t_SLV_LEN : integer := 45;
function uint45_t_to_slv(x : uint45_t) return std_logic_vector;
function slv_to_uint45_t(x : std_logic_vector) return uint45_t;
subtype int45_t is signed(44 downto 0);
constant int45_t_SLV_LEN : integer := 45;
function int45_t_to_slv(x : int45_t) return std_logic_vector;
function slv_to_int45_t(x : std_logic_vector) return int45_t;
subtype uint46_t is unsigned(45 downto 0);
constant uint46_t_SLV_LEN : integer := 46;
function uint46_t_to_slv(x : uint46_t) return std_logic_vector;
function slv_to_uint46_t(x : std_logic_vector) return uint46_t;
subtype int46_t is signed(45 downto 0);
constant int46_t_SLV_LEN : integer := 46;
function int46_t_to_slv(x : int46_t) return std_logic_vector;
function slv_to_int46_t(x : std_logic_vector) return int46_t;
subtype uint47_t is unsigned(46 downto 0);
constant uint47_t_SLV_LEN : integer := 47;
function uint47_t_to_slv(x : uint47_t) return std_logic_vector;
function slv_to_uint47_t(x : std_logic_vector) return uint47_t;
subtype int47_t is signed(46 downto 0);
constant int47_t_SLV_LEN : integer := 47;
function int47_t_to_slv(x : int47_t) return std_logic_vector;
function slv_to_int47_t(x : std_logic_vector) return int47_t;
subtype uint48_t is unsigned(47 downto 0);
constant uint48_t_SLV_LEN : integer := 48;
function uint48_t_to_slv(x : uint48_t) return std_logic_vector;
function slv_to_uint48_t(x : std_logic_vector) return uint48_t;
subtype int48_t is signed(47 downto 0);
constant int48_t_SLV_LEN : integer := 48;
function int48_t_to_slv(x : int48_t) return std_logic_vector;
function slv_to_int48_t(x : std_logic_vector) return int48_t;
subtype uint49_t is unsigned(48 downto 0);
constant uint49_t_SLV_LEN : integer := 49;
function uint49_t_to_slv(x : uint49_t) return std_logic_vector;
function slv_to_uint49_t(x : std_logic_vector) return uint49_t;
subtype int49_t is signed(48 downto 0);
constant int49_t_SLV_LEN : integer := 49;
function int49_t_to_slv(x : int49_t) return std_logic_vector;
function slv_to_int49_t(x : std_logic_vector) return int49_t;
subtype uint50_t is unsigned(49 downto 0);
constant uint50_t_SLV_LEN : integer := 50;
function uint50_t_to_slv(x : uint50_t) return std_logic_vector;
function slv_to_uint50_t(x : std_logic_vector) return uint50_t;
subtype int50_t is signed(49 downto 0);
constant int50_t_SLV_LEN : integer := 50;
function int50_t_to_slv(x : int50_t) return std_logic_vector;
function slv_to_int50_t(x : std_logic_vector) return int50_t;
subtype uint51_t is unsigned(50 downto 0);
constant uint51_t_SLV_LEN : integer := 51;
function uint51_t_to_slv(x : uint51_t) return std_logic_vector;
function slv_to_uint51_t(x : std_logic_vector) return uint51_t;
subtype int51_t is signed(50 downto 0);
constant int51_t_SLV_LEN : integer := 51;
function int51_t_to_slv(x : int51_t) return std_logic_vector;
function slv_to_int51_t(x : std_logic_vector) return int51_t;
subtype uint52_t is unsigned(51 downto 0);
constant uint52_t_SLV_LEN : integer := 52;
function uint52_t_to_slv(x : uint52_t) return std_logic_vector;
function slv_to_uint52_t(x : std_logic_vector) return uint52_t;
subtype int52_t is signed(51 downto 0);
constant int52_t_SLV_LEN : integer := 52;
function int52_t_to_slv(x : int52_t) return std_logic_vector;
function slv_to_int52_t(x : std_logic_vector) return int52_t;
subtype uint53_t is unsigned(52 downto 0);
constant uint53_t_SLV_LEN : integer := 53;
function uint53_t_to_slv(x : uint53_t) return std_logic_vector;
function slv_to_uint53_t(x : std_logic_vector) return uint53_t;
subtype int53_t is signed(52 downto 0);
constant int53_t_SLV_LEN : integer := 53;
function int53_t_to_slv(x : int53_t) return std_logic_vector;
function slv_to_int53_t(x : std_logic_vector) return int53_t;
subtype uint54_t is unsigned(53 downto 0);
constant uint54_t_SLV_LEN : integer := 54;
function uint54_t_to_slv(x : uint54_t) return std_logic_vector;
function slv_to_uint54_t(x : std_logic_vector) return uint54_t;
subtype int54_t is signed(53 downto 0);
constant int54_t_SLV_LEN : integer := 54;
function int54_t_to_slv(x : int54_t) return std_logic_vector;
function slv_to_int54_t(x : std_logic_vector) return int54_t;
subtype uint55_t is unsigned(54 downto 0);
constant uint55_t_SLV_LEN : integer := 55;
function uint55_t_to_slv(x : uint55_t) return std_logic_vector;
function slv_to_uint55_t(x : std_logic_vector) return uint55_t;
subtype int55_t is signed(54 downto 0);
constant int55_t_SLV_LEN : integer := 55;
function int55_t_to_slv(x : int55_t) return std_logic_vector;
function slv_to_int55_t(x : std_logic_vector) return int55_t;
subtype uint56_t is unsigned(55 downto 0);
constant uint56_t_SLV_LEN : integer := 56;
function uint56_t_to_slv(x : uint56_t) return std_logic_vector;
function slv_to_uint56_t(x : std_logic_vector) return uint56_t;
subtype int56_t is signed(55 downto 0);
constant int56_t_SLV_LEN : integer := 56;
function int56_t_to_slv(x : int56_t) return std_logic_vector;
function slv_to_int56_t(x : std_logic_vector) return int56_t;
subtype uint57_t is unsigned(56 downto 0);
constant uint57_t_SLV_LEN : integer := 57;
function uint57_t_to_slv(x : uint57_t) return std_logic_vector;
function slv_to_uint57_t(x : std_logic_vector) return uint57_t;
subtype int57_t is signed(56 downto 0);
constant int57_t_SLV_LEN : integer := 57;
function int57_t_to_slv(x : int57_t) return std_logic_vector;
function slv_to_int57_t(x : std_logic_vector) return int57_t;
subtype uint58_t is unsigned(57 downto 0);
constant uint58_t_SLV_LEN : integer := 58;
function uint58_t_to_slv(x : uint58_t) return std_logic_vector;
function slv_to_uint58_t(x : std_logic_vector) return uint58_t;
subtype int58_t is signed(57 downto 0);
constant int58_t_SLV_LEN : integer := 58;
function int58_t_to_slv(x : int58_t) return std_logic_vector;
function slv_to_int58_t(x : std_logic_vector) return int58_t;
subtype uint59_t is unsigned(58 downto 0);
constant uint59_t_SLV_LEN : integer := 59;
function uint59_t_to_slv(x : uint59_t) return std_logic_vector;
function slv_to_uint59_t(x : std_logic_vector) return uint59_t;
subtype int59_t is signed(58 downto 0);
constant int59_t_SLV_LEN : integer := 59;
function int59_t_to_slv(x : int59_t) return std_logic_vector;
function slv_to_int59_t(x : std_logic_vector) return int59_t;
subtype uint60_t is unsigned(59 downto 0);
constant uint60_t_SLV_LEN : integer := 60;
function uint60_t_to_slv(x : uint60_t) return std_logic_vector;
function slv_to_uint60_t(x : std_logic_vector) return uint60_t;
subtype int60_t is signed(59 downto 0);
constant int60_t_SLV_LEN : integer := 60;
function int60_t_to_slv(x : int60_t) return std_logic_vector;
function slv_to_int60_t(x : std_logic_vector) return int60_t;
subtype uint61_t is unsigned(60 downto 0);
constant uint61_t_SLV_LEN : integer := 61;
function uint61_t_to_slv(x : uint61_t) return std_logic_vector;
function slv_to_uint61_t(x : std_logic_vector) return uint61_t;
subtype int61_t is signed(60 downto 0);
constant int61_t_SLV_LEN : integer := 61;
function int61_t_to_slv(x : int61_t) return std_logic_vector;
function slv_to_int61_t(x : std_logic_vector) return int61_t;
subtype uint62_t is unsigned(61 downto 0);
constant uint62_t_SLV_LEN : integer := 62;
function uint62_t_to_slv(x : uint62_t) return std_logic_vector;
function slv_to_uint62_t(x : std_logic_vector) return uint62_t;
subtype int62_t is signed(61 downto 0);
constant int62_t_SLV_LEN : integer := 62;
function int62_t_to_slv(x : int62_t) return std_logic_vector;
function slv_to_int62_t(x : std_logic_vector) return int62_t;
subtype uint63_t is unsigned(62 downto 0);
constant uint63_t_SLV_LEN : integer := 63;
function uint63_t_to_slv(x : uint63_t) return std_logic_vector;
function slv_to_uint63_t(x : std_logic_vector) return uint63_t;
subtype int63_t is signed(62 downto 0);
constant int63_t_SLV_LEN : integer := 63;
function int63_t_to_slv(x : int63_t) return std_logic_vector;
function slv_to_int63_t(x : std_logic_vector) return int63_t;
subtype uint64_t is unsigned(63 downto 0);
constant uint64_t_SLV_LEN : integer := 64;
function uint64_t_to_slv(x : uint64_t) return std_logic_vector;
function slv_to_uint64_t(x : std_logic_vector) return uint64_t;
subtype int64_t is signed(63 downto 0);
constant int64_t_SLV_LEN : integer := 64;
function int64_t_to_slv(x : int64_t) return std_logic_vector;
function slv_to_int64_t(x : std_logic_vector) return int64_t;
subtype uint65_t is unsigned(64 downto 0);
constant uint65_t_SLV_LEN : integer := 65;
function uint65_t_to_slv(x : uint65_t) return std_logic_vector;
function slv_to_uint65_t(x : std_logic_vector) return uint65_t;
subtype int65_t is signed(64 downto 0);
constant int65_t_SLV_LEN : integer := 65;
function int65_t_to_slv(x : int65_t) return std_logic_vector;
function slv_to_int65_t(x : std_logic_vector) return int65_t;
subtype uint66_t is unsigned(65 downto 0);
constant uint66_t_SLV_LEN : integer := 66;
function uint66_t_to_slv(x : uint66_t) return std_logic_vector;
function slv_to_uint66_t(x : std_logic_vector) return uint66_t;
subtype int66_t is signed(65 downto 0);
constant int66_t_SLV_LEN : integer := 66;
function int66_t_to_slv(x : int66_t) return std_logic_vector;
function slv_to_int66_t(x : std_logic_vector) return int66_t;
subtype uint67_t is unsigned(66 downto 0);
constant uint67_t_SLV_LEN : integer := 67;
function uint67_t_to_slv(x : uint67_t) return std_logic_vector;
function slv_to_uint67_t(x : std_logic_vector) return uint67_t;
subtype int67_t is signed(66 downto 0);
constant int67_t_SLV_LEN : integer := 67;
function int67_t_to_slv(x : int67_t) return std_logic_vector;
function slv_to_int67_t(x : std_logic_vector) return int67_t;
subtype uint68_t is unsigned(67 downto 0);
constant uint68_t_SLV_LEN : integer := 68;
function uint68_t_to_slv(x : uint68_t) return std_logic_vector;
function slv_to_uint68_t(x : std_logic_vector) return uint68_t;
subtype int68_t is signed(67 downto 0);
constant int68_t_SLV_LEN : integer := 68;
function int68_t_to_slv(x : int68_t) return std_logic_vector;
function slv_to_int68_t(x : std_logic_vector) return int68_t;
subtype uint69_t is unsigned(68 downto 0);
constant uint69_t_SLV_LEN : integer := 69;
function uint69_t_to_slv(x : uint69_t) return std_logic_vector;
function slv_to_uint69_t(x : std_logic_vector) return uint69_t;
subtype int69_t is signed(68 downto 0);
constant int69_t_SLV_LEN : integer := 69;
function int69_t_to_slv(x : int69_t) return std_logic_vector;
function slv_to_int69_t(x : std_logic_vector) return int69_t;
subtype uint70_t is unsigned(69 downto 0);
constant uint70_t_SLV_LEN : integer := 70;
function uint70_t_to_slv(x : uint70_t) return std_logic_vector;
function slv_to_uint70_t(x : std_logic_vector) return uint70_t;
subtype int70_t is signed(69 downto 0);
constant int70_t_SLV_LEN : integer := 70;
function int70_t_to_slv(x : int70_t) return std_logic_vector;
function slv_to_int70_t(x : std_logic_vector) return int70_t;
subtype uint71_t is unsigned(70 downto 0);
constant uint71_t_SLV_LEN : integer := 71;
function uint71_t_to_slv(x : uint71_t) return std_logic_vector;
function slv_to_uint71_t(x : std_logic_vector) return uint71_t;
subtype int71_t is signed(70 downto 0);
constant int71_t_SLV_LEN : integer := 71;
function int71_t_to_slv(x : int71_t) return std_logic_vector;
function slv_to_int71_t(x : std_logic_vector) return int71_t;
subtype uint72_t is unsigned(71 downto 0);
constant uint72_t_SLV_LEN : integer := 72;
function uint72_t_to_slv(x : uint72_t) return std_logic_vector;
function slv_to_uint72_t(x : std_logic_vector) return uint72_t;
subtype int72_t is signed(71 downto 0);
constant int72_t_SLV_LEN : integer := 72;
function int72_t_to_slv(x : int72_t) return std_logic_vector;
function slv_to_int72_t(x : std_logic_vector) return int72_t;
subtype uint73_t is unsigned(72 downto 0);
constant uint73_t_SLV_LEN : integer := 73;
function uint73_t_to_slv(x : uint73_t) return std_logic_vector;
function slv_to_uint73_t(x : std_logic_vector) return uint73_t;
subtype int73_t is signed(72 downto 0);
constant int73_t_SLV_LEN : integer := 73;
function int73_t_to_slv(x : int73_t) return std_logic_vector;
function slv_to_int73_t(x : std_logic_vector) return int73_t;
subtype uint74_t is unsigned(73 downto 0);
constant uint74_t_SLV_LEN : integer := 74;
function uint74_t_to_slv(x : uint74_t) return std_logic_vector;
function slv_to_uint74_t(x : std_logic_vector) return uint74_t;
subtype int74_t is signed(73 downto 0);
constant int74_t_SLV_LEN : integer := 74;
function int74_t_to_slv(x : int74_t) return std_logic_vector;
function slv_to_int74_t(x : std_logic_vector) return int74_t;
subtype uint75_t is unsigned(74 downto 0);
constant uint75_t_SLV_LEN : integer := 75;
function uint75_t_to_slv(x : uint75_t) return std_logic_vector;
function slv_to_uint75_t(x : std_logic_vector) return uint75_t;
subtype int75_t is signed(74 downto 0);
constant int75_t_SLV_LEN : integer := 75;
function int75_t_to_slv(x : int75_t) return std_logic_vector;
function slv_to_int75_t(x : std_logic_vector) return int75_t;
subtype uint76_t is unsigned(75 downto 0);
constant uint76_t_SLV_LEN : integer := 76;
function uint76_t_to_slv(x : uint76_t) return std_logic_vector;
function slv_to_uint76_t(x : std_logic_vector) return uint76_t;
subtype int76_t is signed(75 downto 0);
constant int76_t_SLV_LEN : integer := 76;
function int76_t_to_slv(x : int76_t) return std_logic_vector;
function slv_to_int76_t(x : std_logic_vector) return int76_t;
subtype uint77_t is unsigned(76 downto 0);
constant uint77_t_SLV_LEN : integer := 77;
function uint77_t_to_slv(x : uint77_t) return std_logic_vector;
function slv_to_uint77_t(x : std_logic_vector) return uint77_t;
subtype int77_t is signed(76 downto 0);
constant int77_t_SLV_LEN : integer := 77;
function int77_t_to_slv(x : int77_t) return std_logic_vector;
function slv_to_int77_t(x : std_logic_vector) return int77_t;
subtype uint78_t is unsigned(77 downto 0);
constant uint78_t_SLV_LEN : integer := 78;
function uint78_t_to_slv(x : uint78_t) return std_logic_vector;
function slv_to_uint78_t(x : std_logic_vector) return uint78_t;
subtype int78_t is signed(77 downto 0);
constant int78_t_SLV_LEN : integer := 78;
function int78_t_to_slv(x : int78_t) return std_logic_vector;
function slv_to_int78_t(x : std_logic_vector) return int78_t;
subtype uint79_t is unsigned(78 downto 0);
constant uint79_t_SLV_LEN : integer := 79;
function uint79_t_to_slv(x : uint79_t) return std_logic_vector;
function slv_to_uint79_t(x : std_logic_vector) return uint79_t;
subtype int79_t is signed(78 downto 0);
constant int79_t_SLV_LEN : integer := 79;
function int79_t_to_slv(x : int79_t) return std_logic_vector;
function slv_to_int79_t(x : std_logic_vector) return int79_t;
subtype uint80_t is unsigned(79 downto 0);
constant uint80_t_SLV_LEN : integer := 80;
function uint80_t_to_slv(x : uint80_t) return std_logic_vector;
function slv_to_uint80_t(x : std_logic_vector) return uint80_t;
subtype int80_t is signed(79 downto 0);
constant int80_t_SLV_LEN : integer := 80;
function int80_t_to_slv(x : int80_t) return std_logic_vector;
function slv_to_int80_t(x : std_logic_vector) return int80_t;
subtype uint81_t is unsigned(80 downto 0);
constant uint81_t_SLV_LEN : integer := 81;
function uint81_t_to_slv(x : uint81_t) return std_logic_vector;
function slv_to_uint81_t(x : std_logic_vector) return uint81_t;
subtype int81_t is signed(80 downto 0);
constant int81_t_SLV_LEN : integer := 81;
function int81_t_to_slv(x : int81_t) return std_logic_vector;
function slv_to_int81_t(x : std_logic_vector) return int81_t;
subtype uint82_t is unsigned(81 downto 0);
constant uint82_t_SLV_LEN : integer := 82;
function uint82_t_to_slv(x : uint82_t) return std_logic_vector;
function slv_to_uint82_t(x : std_logic_vector) return uint82_t;
subtype int82_t is signed(81 downto 0);
constant int82_t_SLV_LEN : integer := 82;
function int82_t_to_slv(x : int82_t) return std_logic_vector;
function slv_to_int82_t(x : std_logic_vector) return int82_t;
subtype uint83_t is unsigned(82 downto 0);
constant uint83_t_SLV_LEN : integer := 83;
function uint83_t_to_slv(x : uint83_t) return std_logic_vector;
function slv_to_uint83_t(x : std_logic_vector) return uint83_t;
subtype int83_t is signed(82 downto 0);
constant int83_t_SLV_LEN : integer := 83;
function int83_t_to_slv(x : int83_t) return std_logic_vector;
function slv_to_int83_t(x : std_logic_vector) return int83_t;
subtype uint84_t is unsigned(83 downto 0);
constant uint84_t_SLV_LEN : integer := 84;
function uint84_t_to_slv(x : uint84_t) return std_logic_vector;
function slv_to_uint84_t(x : std_logic_vector) return uint84_t;
subtype int84_t is signed(83 downto 0);
constant int84_t_SLV_LEN : integer := 84;
function int84_t_to_slv(x : int84_t) return std_logic_vector;
function slv_to_int84_t(x : std_logic_vector) return int84_t;
subtype uint85_t is unsigned(84 downto 0);
constant uint85_t_SLV_LEN : integer := 85;
function uint85_t_to_slv(x : uint85_t) return std_logic_vector;
function slv_to_uint85_t(x : std_logic_vector) return uint85_t;
subtype int85_t is signed(84 downto 0);
constant int85_t_SLV_LEN : integer := 85;
function int85_t_to_slv(x : int85_t) return std_logic_vector;
function slv_to_int85_t(x : std_logic_vector) return int85_t;
subtype uint86_t is unsigned(85 downto 0);
constant uint86_t_SLV_LEN : integer := 86;
function uint86_t_to_slv(x : uint86_t) return std_logic_vector;
function slv_to_uint86_t(x : std_logic_vector) return uint86_t;
subtype int86_t is signed(85 downto 0);
constant int86_t_SLV_LEN : integer := 86;
function int86_t_to_slv(x : int86_t) return std_logic_vector;
function slv_to_int86_t(x : std_logic_vector) return int86_t;
subtype uint87_t is unsigned(86 downto 0);
constant uint87_t_SLV_LEN : integer := 87;
function uint87_t_to_slv(x : uint87_t) return std_logic_vector;
function slv_to_uint87_t(x : std_logic_vector) return uint87_t;
subtype int87_t is signed(86 downto 0);
constant int87_t_SLV_LEN : integer := 87;
function int87_t_to_slv(x : int87_t) return std_logic_vector;
function slv_to_int87_t(x : std_logic_vector) return int87_t;
subtype uint88_t is unsigned(87 downto 0);
constant uint88_t_SLV_LEN : integer := 88;
function uint88_t_to_slv(x : uint88_t) return std_logic_vector;
function slv_to_uint88_t(x : std_logic_vector) return uint88_t;
subtype int88_t is signed(87 downto 0);
constant int88_t_SLV_LEN : integer := 88;
function int88_t_to_slv(x : int88_t) return std_logic_vector;
function slv_to_int88_t(x : std_logic_vector) return int88_t;
subtype uint89_t is unsigned(88 downto 0);
constant uint89_t_SLV_LEN : integer := 89;
function uint89_t_to_slv(x : uint89_t) return std_logic_vector;
function slv_to_uint89_t(x : std_logic_vector) return uint89_t;
subtype int89_t is signed(88 downto 0);
constant int89_t_SLV_LEN : integer := 89;
function int89_t_to_slv(x : int89_t) return std_logic_vector;
function slv_to_int89_t(x : std_logic_vector) return int89_t;
subtype uint90_t is unsigned(89 downto 0);
constant uint90_t_SLV_LEN : integer := 90;
function uint90_t_to_slv(x : uint90_t) return std_logic_vector;
function slv_to_uint90_t(x : std_logic_vector) return uint90_t;
subtype int90_t is signed(89 downto 0);
constant int90_t_SLV_LEN : integer := 90;
function int90_t_to_slv(x : int90_t) return std_logic_vector;
function slv_to_int90_t(x : std_logic_vector) return int90_t;
subtype uint91_t is unsigned(90 downto 0);
constant uint91_t_SLV_LEN : integer := 91;
function uint91_t_to_slv(x : uint91_t) return std_logic_vector;
function slv_to_uint91_t(x : std_logic_vector) return uint91_t;
subtype int91_t is signed(90 downto 0);
constant int91_t_SLV_LEN : integer := 91;
function int91_t_to_slv(x : int91_t) return std_logic_vector;
function slv_to_int91_t(x : std_logic_vector) return int91_t;
subtype uint92_t is unsigned(91 downto 0);
constant uint92_t_SLV_LEN : integer := 92;
function uint92_t_to_slv(x : uint92_t) return std_logic_vector;
function slv_to_uint92_t(x : std_logic_vector) return uint92_t;
subtype int92_t is signed(91 downto 0);
constant int92_t_SLV_LEN : integer := 92;
function int92_t_to_slv(x : int92_t) return std_logic_vector;
function slv_to_int92_t(x : std_logic_vector) return int92_t;
subtype uint93_t is unsigned(92 downto 0);
constant uint93_t_SLV_LEN : integer := 93;
function uint93_t_to_slv(x : uint93_t) return std_logic_vector;
function slv_to_uint93_t(x : std_logic_vector) return uint93_t;
subtype int93_t is signed(92 downto 0);
constant int93_t_SLV_LEN : integer := 93;
function int93_t_to_slv(x : int93_t) return std_logic_vector;
function slv_to_int93_t(x : std_logic_vector) return int93_t;
subtype uint94_t is unsigned(93 downto 0);
constant uint94_t_SLV_LEN : integer := 94;
function uint94_t_to_slv(x : uint94_t) return std_logic_vector;
function slv_to_uint94_t(x : std_logic_vector) return uint94_t;
subtype int94_t is signed(93 downto 0);
constant int94_t_SLV_LEN : integer := 94;
function int94_t_to_slv(x : int94_t) return std_logic_vector;
function slv_to_int94_t(x : std_logic_vector) return int94_t;
subtype uint95_t is unsigned(94 downto 0);
constant uint95_t_SLV_LEN : integer := 95;
function uint95_t_to_slv(x : uint95_t) return std_logic_vector;
function slv_to_uint95_t(x : std_logic_vector) return uint95_t;
subtype int95_t is signed(94 downto 0);
constant int95_t_SLV_LEN : integer := 95;
function int95_t_to_slv(x : int95_t) return std_logic_vector;
function slv_to_int95_t(x : std_logic_vector) return int95_t;
subtype uint96_t is unsigned(95 downto 0);
constant uint96_t_SLV_LEN : integer := 96;
function uint96_t_to_slv(x : uint96_t) return std_logic_vector;
function slv_to_uint96_t(x : std_logic_vector) return uint96_t;
subtype int96_t is signed(95 downto 0);
constant int96_t_SLV_LEN : integer := 96;
function int96_t_to_slv(x : int96_t) return std_logic_vector;
function slv_to_int96_t(x : std_logic_vector) return int96_t;
subtype uint97_t is unsigned(96 downto 0);
constant uint97_t_SLV_LEN : integer := 97;
function uint97_t_to_slv(x : uint97_t) return std_logic_vector;
function slv_to_uint97_t(x : std_logic_vector) return uint97_t;
subtype int97_t is signed(96 downto 0);
constant int97_t_SLV_LEN : integer := 97;
function int97_t_to_slv(x : int97_t) return std_logic_vector;
function slv_to_int97_t(x : std_logic_vector) return int97_t;
subtype uint98_t is unsigned(97 downto 0);
constant uint98_t_SLV_LEN : integer := 98;
function uint98_t_to_slv(x : uint98_t) return std_logic_vector;
function slv_to_uint98_t(x : std_logic_vector) return uint98_t;
subtype int98_t is signed(97 downto 0);
constant int98_t_SLV_LEN : integer := 98;
function int98_t_to_slv(x : int98_t) return std_logic_vector;
function slv_to_int98_t(x : std_logic_vector) return int98_t;
subtype uint99_t is unsigned(98 downto 0);
constant uint99_t_SLV_LEN : integer := 99;
function uint99_t_to_slv(x : uint99_t) return std_logic_vector;
function slv_to_uint99_t(x : std_logic_vector) return uint99_t;
subtype int99_t is signed(98 downto 0);
constant int99_t_SLV_LEN : integer := 99;
function int99_t_to_slv(x : int99_t) return std_logic_vector;
function slv_to_int99_t(x : std_logic_vector) return int99_t;
subtype uint100_t is unsigned(99 downto 0);
constant uint100_t_SLV_LEN : integer := 100;
function uint100_t_to_slv(x : uint100_t) return std_logic_vector;
function slv_to_uint100_t(x : std_logic_vector) return uint100_t;
subtype int100_t is signed(99 downto 0);
constant int100_t_SLV_LEN : integer := 100;
function int100_t_to_slv(x : int100_t) return std_logic_vector;
function slv_to_int100_t(x : std_logic_vector) return int100_t;
subtype uint101_t is unsigned(100 downto 0);
constant uint101_t_SLV_LEN : integer := 101;
function uint101_t_to_slv(x : uint101_t) return std_logic_vector;
function slv_to_uint101_t(x : std_logic_vector) return uint101_t;
subtype int101_t is signed(100 downto 0);
constant int101_t_SLV_LEN : integer := 101;
function int101_t_to_slv(x : int101_t) return std_logic_vector;
function slv_to_int101_t(x : std_logic_vector) return int101_t;
subtype uint102_t is unsigned(101 downto 0);
constant uint102_t_SLV_LEN : integer := 102;
function uint102_t_to_slv(x : uint102_t) return std_logic_vector;
function slv_to_uint102_t(x : std_logic_vector) return uint102_t;
subtype int102_t is signed(101 downto 0);
constant int102_t_SLV_LEN : integer := 102;
function int102_t_to_slv(x : int102_t) return std_logic_vector;
function slv_to_int102_t(x : std_logic_vector) return int102_t;
subtype uint103_t is unsigned(102 downto 0);
constant uint103_t_SLV_LEN : integer := 103;
function uint103_t_to_slv(x : uint103_t) return std_logic_vector;
function slv_to_uint103_t(x : std_logic_vector) return uint103_t;
subtype int103_t is signed(102 downto 0);
constant int103_t_SLV_LEN : integer := 103;
function int103_t_to_slv(x : int103_t) return std_logic_vector;
function slv_to_int103_t(x : std_logic_vector) return int103_t;
subtype uint104_t is unsigned(103 downto 0);
constant uint104_t_SLV_LEN : integer := 104;
function uint104_t_to_slv(x : uint104_t) return std_logic_vector;
function slv_to_uint104_t(x : std_logic_vector) return uint104_t;
subtype int104_t is signed(103 downto 0);
constant int104_t_SLV_LEN : integer := 104;
function int104_t_to_slv(x : int104_t) return std_logic_vector;
function slv_to_int104_t(x : std_logic_vector) return int104_t;
subtype uint105_t is unsigned(104 downto 0);
constant uint105_t_SLV_LEN : integer := 105;
function uint105_t_to_slv(x : uint105_t) return std_logic_vector;
function slv_to_uint105_t(x : std_logic_vector) return uint105_t;
subtype int105_t is signed(104 downto 0);
constant int105_t_SLV_LEN : integer := 105;
function int105_t_to_slv(x : int105_t) return std_logic_vector;
function slv_to_int105_t(x : std_logic_vector) return int105_t;
subtype uint106_t is unsigned(105 downto 0);
constant uint106_t_SLV_LEN : integer := 106;
function uint106_t_to_slv(x : uint106_t) return std_logic_vector;
function slv_to_uint106_t(x : std_logic_vector) return uint106_t;
subtype int106_t is signed(105 downto 0);
constant int106_t_SLV_LEN : integer := 106;
function int106_t_to_slv(x : int106_t) return std_logic_vector;
function slv_to_int106_t(x : std_logic_vector) return int106_t;
subtype uint107_t is unsigned(106 downto 0);
constant uint107_t_SLV_LEN : integer := 107;
function uint107_t_to_slv(x : uint107_t) return std_logic_vector;
function slv_to_uint107_t(x : std_logic_vector) return uint107_t;
subtype int107_t is signed(106 downto 0);
constant int107_t_SLV_LEN : integer := 107;
function int107_t_to_slv(x : int107_t) return std_logic_vector;
function slv_to_int107_t(x : std_logic_vector) return int107_t;
subtype uint108_t is unsigned(107 downto 0);
constant uint108_t_SLV_LEN : integer := 108;
function uint108_t_to_slv(x : uint108_t) return std_logic_vector;
function slv_to_uint108_t(x : std_logic_vector) return uint108_t;
subtype int108_t is signed(107 downto 0);
constant int108_t_SLV_LEN : integer := 108;
function int108_t_to_slv(x : int108_t) return std_logic_vector;
function slv_to_int108_t(x : std_logic_vector) return int108_t;
subtype uint109_t is unsigned(108 downto 0);
constant uint109_t_SLV_LEN : integer := 109;
function uint109_t_to_slv(x : uint109_t) return std_logic_vector;
function slv_to_uint109_t(x : std_logic_vector) return uint109_t;
subtype int109_t is signed(108 downto 0);
constant int109_t_SLV_LEN : integer := 109;
function int109_t_to_slv(x : int109_t) return std_logic_vector;
function slv_to_int109_t(x : std_logic_vector) return int109_t;
subtype uint110_t is unsigned(109 downto 0);
constant uint110_t_SLV_LEN : integer := 110;
function uint110_t_to_slv(x : uint110_t) return std_logic_vector;
function slv_to_uint110_t(x : std_logic_vector) return uint110_t;
subtype int110_t is signed(109 downto 0);
constant int110_t_SLV_LEN : integer := 110;
function int110_t_to_slv(x : int110_t) return std_logic_vector;
function slv_to_int110_t(x : std_logic_vector) return int110_t;
subtype uint111_t is unsigned(110 downto 0);
constant uint111_t_SLV_LEN : integer := 111;
function uint111_t_to_slv(x : uint111_t) return std_logic_vector;
function slv_to_uint111_t(x : std_logic_vector) return uint111_t;
subtype int111_t is signed(110 downto 0);
constant int111_t_SLV_LEN : integer := 111;
function int111_t_to_slv(x : int111_t) return std_logic_vector;
function slv_to_int111_t(x : std_logic_vector) return int111_t;
subtype uint112_t is unsigned(111 downto 0);
constant uint112_t_SLV_LEN : integer := 112;
function uint112_t_to_slv(x : uint112_t) return std_logic_vector;
function slv_to_uint112_t(x : std_logic_vector) return uint112_t;
subtype int112_t is signed(111 downto 0);
constant int112_t_SLV_LEN : integer := 112;
function int112_t_to_slv(x : int112_t) return std_logic_vector;
function slv_to_int112_t(x : std_logic_vector) return int112_t;
subtype uint113_t is unsigned(112 downto 0);
constant uint113_t_SLV_LEN : integer := 113;
function uint113_t_to_slv(x : uint113_t) return std_logic_vector;
function slv_to_uint113_t(x : std_logic_vector) return uint113_t;
subtype int113_t is signed(112 downto 0);
constant int113_t_SLV_LEN : integer := 113;
function int113_t_to_slv(x : int113_t) return std_logic_vector;
function slv_to_int113_t(x : std_logic_vector) return int113_t;
subtype uint114_t is unsigned(113 downto 0);
constant uint114_t_SLV_LEN : integer := 114;
function uint114_t_to_slv(x : uint114_t) return std_logic_vector;
function slv_to_uint114_t(x : std_logic_vector) return uint114_t;
subtype int114_t is signed(113 downto 0);
constant int114_t_SLV_LEN : integer := 114;
function int114_t_to_slv(x : int114_t) return std_logic_vector;
function slv_to_int114_t(x : std_logic_vector) return int114_t;
subtype uint115_t is unsigned(114 downto 0);
constant uint115_t_SLV_LEN : integer := 115;
function uint115_t_to_slv(x : uint115_t) return std_logic_vector;
function slv_to_uint115_t(x : std_logic_vector) return uint115_t;
subtype int115_t is signed(114 downto 0);
constant int115_t_SLV_LEN : integer := 115;
function int115_t_to_slv(x : int115_t) return std_logic_vector;
function slv_to_int115_t(x : std_logic_vector) return int115_t;
subtype uint116_t is unsigned(115 downto 0);
constant uint116_t_SLV_LEN : integer := 116;
function uint116_t_to_slv(x : uint116_t) return std_logic_vector;
function slv_to_uint116_t(x : std_logic_vector) return uint116_t;
subtype int116_t is signed(115 downto 0);
constant int116_t_SLV_LEN : integer := 116;
function int116_t_to_slv(x : int116_t) return std_logic_vector;
function slv_to_int116_t(x : std_logic_vector) return int116_t;
subtype uint117_t is unsigned(116 downto 0);
constant uint117_t_SLV_LEN : integer := 117;
function uint117_t_to_slv(x : uint117_t) return std_logic_vector;
function slv_to_uint117_t(x : std_logic_vector) return uint117_t;
subtype int117_t is signed(116 downto 0);
constant int117_t_SLV_LEN : integer := 117;
function int117_t_to_slv(x : int117_t) return std_logic_vector;
function slv_to_int117_t(x : std_logic_vector) return int117_t;
subtype uint118_t is unsigned(117 downto 0);
constant uint118_t_SLV_LEN : integer := 118;
function uint118_t_to_slv(x : uint118_t) return std_logic_vector;
function slv_to_uint118_t(x : std_logic_vector) return uint118_t;
subtype int118_t is signed(117 downto 0);
constant int118_t_SLV_LEN : integer := 118;
function int118_t_to_slv(x : int118_t) return std_logic_vector;
function slv_to_int118_t(x : std_logic_vector) return int118_t;
subtype uint119_t is unsigned(118 downto 0);
constant uint119_t_SLV_LEN : integer := 119;
function uint119_t_to_slv(x : uint119_t) return std_logic_vector;
function slv_to_uint119_t(x : std_logic_vector) return uint119_t;
subtype int119_t is signed(118 downto 0);
constant int119_t_SLV_LEN : integer := 119;
function int119_t_to_slv(x : int119_t) return std_logic_vector;
function slv_to_int119_t(x : std_logic_vector) return int119_t;
subtype uint120_t is unsigned(119 downto 0);
constant uint120_t_SLV_LEN : integer := 120;
function uint120_t_to_slv(x : uint120_t) return std_logic_vector;
function slv_to_uint120_t(x : std_logic_vector) return uint120_t;
subtype int120_t is signed(119 downto 0);
constant int120_t_SLV_LEN : integer := 120;
function int120_t_to_slv(x : int120_t) return std_logic_vector;
function slv_to_int120_t(x : std_logic_vector) return int120_t;
subtype uint121_t is unsigned(120 downto 0);
constant uint121_t_SLV_LEN : integer := 121;
function uint121_t_to_slv(x : uint121_t) return std_logic_vector;
function slv_to_uint121_t(x : std_logic_vector) return uint121_t;
subtype int121_t is signed(120 downto 0);
constant int121_t_SLV_LEN : integer := 121;
function int121_t_to_slv(x : int121_t) return std_logic_vector;
function slv_to_int121_t(x : std_logic_vector) return int121_t;
subtype uint122_t is unsigned(121 downto 0);
constant uint122_t_SLV_LEN : integer := 122;
function uint122_t_to_slv(x : uint122_t) return std_logic_vector;
function slv_to_uint122_t(x : std_logic_vector) return uint122_t;
subtype int122_t is signed(121 downto 0);
constant int122_t_SLV_LEN : integer := 122;
function int122_t_to_slv(x : int122_t) return std_logic_vector;
function slv_to_int122_t(x : std_logic_vector) return int122_t;
subtype uint123_t is unsigned(122 downto 0);
constant uint123_t_SLV_LEN : integer := 123;
function uint123_t_to_slv(x : uint123_t) return std_logic_vector;
function slv_to_uint123_t(x : std_logic_vector) return uint123_t;
subtype int123_t is signed(122 downto 0);
constant int123_t_SLV_LEN : integer := 123;
function int123_t_to_slv(x : int123_t) return std_logic_vector;
function slv_to_int123_t(x : std_logic_vector) return int123_t;
subtype uint124_t is unsigned(123 downto 0);
constant uint124_t_SLV_LEN : integer := 124;
function uint124_t_to_slv(x : uint124_t) return std_logic_vector;
function slv_to_uint124_t(x : std_logic_vector) return uint124_t;
subtype int124_t is signed(123 downto 0);
constant int124_t_SLV_LEN : integer := 124;
function int124_t_to_slv(x : int124_t) return std_logic_vector;
function slv_to_int124_t(x : std_logic_vector) return int124_t;
subtype uint125_t is unsigned(124 downto 0);
constant uint125_t_SLV_LEN : integer := 125;
function uint125_t_to_slv(x : uint125_t) return std_logic_vector;
function slv_to_uint125_t(x : std_logic_vector) return uint125_t;
subtype int125_t is signed(124 downto 0);
constant int125_t_SLV_LEN : integer := 125;
function int125_t_to_slv(x : int125_t) return std_logic_vector;
function slv_to_int125_t(x : std_logic_vector) return int125_t;
subtype uint126_t is unsigned(125 downto 0);
constant uint126_t_SLV_LEN : integer := 126;
function uint126_t_to_slv(x : uint126_t) return std_logic_vector;
function slv_to_uint126_t(x : std_logic_vector) return uint126_t;
subtype int126_t is signed(125 downto 0);
constant int126_t_SLV_LEN : integer := 126;
function int126_t_to_slv(x : int126_t) return std_logic_vector;
function slv_to_int126_t(x : std_logic_vector) return int126_t;
subtype uint127_t is unsigned(126 downto 0);
constant uint127_t_SLV_LEN : integer := 127;
function uint127_t_to_slv(x : uint127_t) return std_logic_vector;
function slv_to_uint127_t(x : std_logic_vector) return uint127_t;
subtype int127_t is signed(126 downto 0);
constant int127_t_SLV_LEN : integer := 127;
function int127_t_to_slv(x : int127_t) return std_logic_vector;
function slv_to_int127_t(x : std_logic_vector) return int127_t;
subtype uint128_t is unsigned(127 downto 0);
constant uint128_t_SLV_LEN : integer := 128;
function uint128_t_to_slv(x : uint128_t) return std_logic_vector;
function slv_to_uint128_t(x : std_logic_vector) return uint128_t;
subtype int128_t is signed(127 downto 0);
constant int128_t_SLV_LEN : integer := 128;
function int128_t_to_slv(x : int128_t) return std_logic_vector;
function slv_to_int128_t(x : std_logic_vector) return int128_t;
subtype uint129_t is unsigned(128 downto 0);
constant uint129_t_SLV_LEN : integer := 129;
function uint129_t_to_slv(x : uint129_t) return std_logic_vector;
function slv_to_uint129_t(x : std_logic_vector) return uint129_t;
subtype int129_t is signed(128 downto 0);
constant int129_t_SLV_LEN : integer := 129;
function int129_t_to_slv(x : int129_t) return std_logic_vector;
function slv_to_int129_t(x : std_logic_vector) return int129_t;
subtype uint130_t is unsigned(129 downto 0);
constant uint130_t_SLV_LEN : integer := 130;
function uint130_t_to_slv(x : uint130_t) return std_logic_vector;
function slv_to_uint130_t(x : std_logic_vector) return uint130_t;
subtype int130_t is signed(129 downto 0);
constant int130_t_SLV_LEN : integer := 130;
function int130_t_to_slv(x : int130_t) return std_logic_vector;
function slv_to_int130_t(x : std_logic_vector) return int130_t;
subtype uint131_t is unsigned(130 downto 0);
constant uint131_t_SLV_LEN : integer := 131;
function uint131_t_to_slv(x : uint131_t) return std_logic_vector;
function slv_to_uint131_t(x : std_logic_vector) return uint131_t;
subtype int131_t is signed(130 downto 0);
constant int131_t_SLV_LEN : integer := 131;
function int131_t_to_slv(x : int131_t) return std_logic_vector;
function slv_to_int131_t(x : std_logic_vector) return int131_t;
subtype uint132_t is unsigned(131 downto 0);
constant uint132_t_SLV_LEN : integer := 132;
function uint132_t_to_slv(x : uint132_t) return std_logic_vector;
function slv_to_uint132_t(x : std_logic_vector) return uint132_t;
subtype int132_t is signed(131 downto 0);
constant int132_t_SLV_LEN : integer := 132;
function int132_t_to_slv(x : int132_t) return std_logic_vector;
function slv_to_int132_t(x : std_logic_vector) return int132_t;
subtype uint133_t is unsigned(132 downto 0);
constant uint133_t_SLV_LEN : integer := 133;
function uint133_t_to_slv(x : uint133_t) return std_logic_vector;
function slv_to_uint133_t(x : std_logic_vector) return uint133_t;
subtype int133_t is signed(132 downto 0);
constant int133_t_SLV_LEN : integer := 133;
function int133_t_to_slv(x : int133_t) return std_logic_vector;
function slv_to_int133_t(x : std_logic_vector) return int133_t;
subtype uint134_t is unsigned(133 downto 0);
constant uint134_t_SLV_LEN : integer := 134;
function uint134_t_to_slv(x : uint134_t) return std_logic_vector;
function slv_to_uint134_t(x : std_logic_vector) return uint134_t;
subtype int134_t is signed(133 downto 0);
constant int134_t_SLV_LEN : integer := 134;
function int134_t_to_slv(x : int134_t) return std_logic_vector;
function slv_to_int134_t(x : std_logic_vector) return int134_t;
subtype uint135_t is unsigned(134 downto 0);
constant uint135_t_SLV_LEN : integer := 135;
function uint135_t_to_slv(x : uint135_t) return std_logic_vector;
function slv_to_uint135_t(x : std_logic_vector) return uint135_t;
subtype int135_t is signed(134 downto 0);
constant int135_t_SLV_LEN : integer := 135;
function int135_t_to_slv(x : int135_t) return std_logic_vector;
function slv_to_int135_t(x : std_logic_vector) return int135_t;
subtype uint136_t is unsigned(135 downto 0);
constant uint136_t_SLV_LEN : integer := 136;
function uint136_t_to_slv(x : uint136_t) return std_logic_vector;
function slv_to_uint136_t(x : std_logic_vector) return uint136_t;
subtype int136_t is signed(135 downto 0);
constant int136_t_SLV_LEN : integer := 136;
function int136_t_to_slv(x : int136_t) return std_logic_vector;
function slv_to_int136_t(x : std_logic_vector) return int136_t;
subtype uint137_t is unsigned(136 downto 0);
constant uint137_t_SLV_LEN : integer := 137;
function uint137_t_to_slv(x : uint137_t) return std_logic_vector;
function slv_to_uint137_t(x : std_logic_vector) return uint137_t;
subtype int137_t is signed(136 downto 0);
constant int137_t_SLV_LEN : integer := 137;
function int137_t_to_slv(x : int137_t) return std_logic_vector;
function slv_to_int137_t(x : std_logic_vector) return int137_t;
subtype uint138_t is unsigned(137 downto 0);
constant uint138_t_SLV_LEN : integer := 138;
function uint138_t_to_slv(x : uint138_t) return std_logic_vector;
function slv_to_uint138_t(x : std_logic_vector) return uint138_t;
subtype int138_t is signed(137 downto 0);
constant int138_t_SLV_LEN : integer := 138;
function int138_t_to_slv(x : int138_t) return std_logic_vector;
function slv_to_int138_t(x : std_logic_vector) return int138_t;
subtype uint139_t is unsigned(138 downto 0);
constant uint139_t_SLV_LEN : integer := 139;
function uint139_t_to_slv(x : uint139_t) return std_logic_vector;
function slv_to_uint139_t(x : std_logic_vector) return uint139_t;
subtype int139_t is signed(138 downto 0);
constant int139_t_SLV_LEN : integer := 139;
function int139_t_to_slv(x : int139_t) return std_logic_vector;
function slv_to_int139_t(x : std_logic_vector) return int139_t;
subtype uint140_t is unsigned(139 downto 0);
constant uint140_t_SLV_LEN : integer := 140;
function uint140_t_to_slv(x : uint140_t) return std_logic_vector;
function slv_to_uint140_t(x : std_logic_vector) return uint140_t;
subtype int140_t is signed(139 downto 0);
constant int140_t_SLV_LEN : integer := 140;
function int140_t_to_slv(x : int140_t) return std_logic_vector;
function slv_to_int140_t(x : std_logic_vector) return int140_t;
subtype uint141_t is unsigned(140 downto 0);
constant uint141_t_SLV_LEN : integer := 141;
function uint141_t_to_slv(x : uint141_t) return std_logic_vector;
function slv_to_uint141_t(x : std_logic_vector) return uint141_t;
subtype int141_t is signed(140 downto 0);
constant int141_t_SLV_LEN : integer := 141;
function int141_t_to_slv(x : int141_t) return std_logic_vector;
function slv_to_int141_t(x : std_logic_vector) return int141_t;
subtype uint142_t is unsigned(141 downto 0);
constant uint142_t_SLV_LEN : integer := 142;
function uint142_t_to_slv(x : uint142_t) return std_logic_vector;
function slv_to_uint142_t(x : std_logic_vector) return uint142_t;
subtype int142_t is signed(141 downto 0);
constant int142_t_SLV_LEN : integer := 142;
function int142_t_to_slv(x : int142_t) return std_logic_vector;
function slv_to_int142_t(x : std_logic_vector) return int142_t;
subtype uint143_t is unsigned(142 downto 0);
constant uint143_t_SLV_LEN : integer := 143;
function uint143_t_to_slv(x : uint143_t) return std_logic_vector;
function slv_to_uint143_t(x : std_logic_vector) return uint143_t;
subtype int143_t is signed(142 downto 0);
constant int143_t_SLV_LEN : integer := 143;
function int143_t_to_slv(x : int143_t) return std_logic_vector;
function slv_to_int143_t(x : std_logic_vector) return int143_t;
subtype uint144_t is unsigned(143 downto 0);
constant uint144_t_SLV_LEN : integer := 144;
function uint144_t_to_slv(x : uint144_t) return std_logic_vector;
function slv_to_uint144_t(x : std_logic_vector) return uint144_t;
subtype int144_t is signed(143 downto 0);
constant int144_t_SLV_LEN : integer := 144;
function int144_t_to_slv(x : int144_t) return std_logic_vector;
function slv_to_int144_t(x : std_logic_vector) return int144_t;
subtype uint145_t is unsigned(144 downto 0);
constant uint145_t_SLV_LEN : integer := 145;
function uint145_t_to_slv(x : uint145_t) return std_logic_vector;
function slv_to_uint145_t(x : std_logic_vector) return uint145_t;
subtype int145_t is signed(144 downto 0);
constant int145_t_SLV_LEN : integer := 145;
function int145_t_to_slv(x : int145_t) return std_logic_vector;
function slv_to_int145_t(x : std_logic_vector) return int145_t;
subtype uint146_t is unsigned(145 downto 0);
constant uint146_t_SLV_LEN : integer := 146;
function uint146_t_to_slv(x : uint146_t) return std_logic_vector;
function slv_to_uint146_t(x : std_logic_vector) return uint146_t;
subtype int146_t is signed(145 downto 0);
constant int146_t_SLV_LEN : integer := 146;
function int146_t_to_slv(x : int146_t) return std_logic_vector;
function slv_to_int146_t(x : std_logic_vector) return int146_t;
subtype uint147_t is unsigned(146 downto 0);
constant uint147_t_SLV_LEN : integer := 147;
function uint147_t_to_slv(x : uint147_t) return std_logic_vector;
function slv_to_uint147_t(x : std_logic_vector) return uint147_t;
subtype int147_t is signed(146 downto 0);
constant int147_t_SLV_LEN : integer := 147;
function int147_t_to_slv(x : int147_t) return std_logic_vector;
function slv_to_int147_t(x : std_logic_vector) return int147_t;
subtype uint148_t is unsigned(147 downto 0);
constant uint148_t_SLV_LEN : integer := 148;
function uint148_t_to_slv(x : uint148_t) return std_logic_vector;
function slv_to_uint148_t(x : std_logic_vector) return uint148_t;
subtype int148_t is signed(147 downto 0);
constant int148_t_SLV_LEN : integer := 148;
function int148_t_to_slv(x : int148_t) return std_logic_vector;
function slv_to_int148_t(x : std_logic_vector) return int148_t;
subtype uint149_t is unsigned(148 downto 0);
constant uint149_t_SLV_LEN : integer := 149;
function uint149_t_to_slv(x : uint149_t) return std_logic_vector;
function slv_to_uint149_t(x : std_logic_vector) return uint149_t;
subtype int149_t is signed(148 downto 0);
constant int149_t_SLV_LEN : integer := 149;
function int149_t_to_slv(x : int149_t) return std_logic_vector;
function slv_to_int149_t(x : std_logic_vector) return int149_t;
subtype uint150_t is unsigned(149 downto 0);
constant uint150_t_SLV_LEN : integer := 150;
function uint150_t_to_slv(x : uint150_t) return std_logic_vector;
function slv_to_uint150_t(x : std_logic_vector) return uint150_t;
subtype int150_t is signed(149 downto 0);
constant int150_t_SLV_LEN : integer := 150;
function int150_t_to_slv(x : int150_t) return std_logic_vector;
function slv_to_int150_t(x : std_logic_vector) return int150_t;
subtype uint151_t is unsigned(150 downto 0);
constant uint151_t_SLV_LEN : integer := 151;
function uint151_t_to_slv(x : uint151_t) return std_logic_vector;
function slv_to_uint151_t(x : std_logic_vector) return uint151_t;
subtype int151_t is signed(150 downto 0);
constant int151_t_SLV_LEN : integer := 151;
function int151_t_to_slv(x : int151_t) return std_logic_vector;
function slv_to_int151_t(x : std_logic_vector) return int151_t;
subtype uint152_t is unsigned(151 downto 0);
constant uint152_t_SLV_LEN : integer := 152;
function uint152_t_to_slv(x : uint152_t) return std_logic_vector;
function slv_to_uint152_t(x : std_logic_vector) return uint152_t;
subtype int152_t is signed(151 downto 0);
constant int152_t_SLV_LEN : integer := 152;
function int152_t_to_slv(x : int152_t) return std_logic_vector;
function slv_to_int152_t(x : std_logic_vector) return int152_t;
subtype uint153_t is unsigned(152 downto 0);
constant uint153_t_SLV_LEN : integer := 153;
function uint153_t_to_slv(x : uint153_t) return std_logic_vector;
function slv_to_uint153_t(x : std_logic_vector) return uint153_t;
subtype int153_t is signed(152 downto 0);
constant int153_t_SLV_LEN : integer := 153;
function int153_t_to_slv(x : int153_t) return std_logic_vector;
function slv_to_int153_t(x : std_logic_vector) return int153_t;
subtype uint154_t is unsigned(153 downto 0);
constant uint154_t_SLV_LEN : integer := 154;
function uint154_t_to_slv(x : uint154_t) return std_logic_vector;
function slv_to_uint154_t(x : std_logic_vector) return uint154_t;
subtype int154_t is signed(153 downto 0);
constant int154_t_SLV_LEN : integer := 154;
function int154_t_to_slv(x : int154_t) return std_logic_vector;
function slv_to_int154_t(x : std_logic_vector) return int154_t;
subtype uint155_t is unsigned(154 downto 0);
constant uint155_t_SLV_LEN : integer := 155;
function uint155_t_to_slv(x : uint155_t) return std_logic_vector;
function slv_to_uint155_t(x : std_logic_vector) return uint155_t;
subtype int155_t is signed(154 downto 0);
constant int155_t_SLV_LEN : integer := 155;
function int155_t_to_slv(x : int155_t) return std_logic_vector;
function slv_to_int155_t(x : std_logic_vector) return int155_t;
subtype uint156_t is unsigned(155 downto 0);
constant uint156_t_SLV_LEN : integer := 156;
function uint156_t_to_slv(x : uint156_t) return std_logic_vector;
function slv_to_uint156_t(x : std_logic_vector) return uint156_t;
subtype int156_t is signed(155 downto 0);
constant int156_t_SLV_LEN : integer := 156;
function int156_t_to_slv(x : int156_t) return std_logic_vector;
function slv_to_int156_t(x : std_logic_vector) return int156_t;
subtype uint157_t is unsigned(156 downto 0);
constant uint157_t_SLV_LEN : integer := 157;
function uint157_t_to_slv(x : uint157_t) return std_logic_vector;
function slv_to_uint157_t(x : std_logic_vector) return uint157_t;
subtype int157_t is signed(156 downto 0);
constant int157_t_SLV_LEN : integer := 157;
function int157_t_to_slv(x : int157_t) return std_logic_vector;
function slv_to_int157_t(x : std_logic_vector) return int157_t;
subtype uint158_t is unsigned(157 downto 0);
constant uint158_t_SLV_LEN : integer := 158;
function uint158_t_to_slv(x : uint158_t) return std_logic_vector;
function slv_to_uint158_t(x : std_logic_vector) return uint158_t;
subtype int158_t is signed(157 downto 0);
constant int158_t_SLV_LEN : integer := 158;
function int158_t_to_slv(x : int158_t) return std_logic_vector;
function slv_to_int158_t(x : std_logic_vector) return int158_t;
subtype uint159_t is unsigned(158 downto 0);
constant uint159_t_SLV_LEN : integer := 159;
function uint159_t_to_slv(x : uint159_t) return std_logic_vector;
function slv_to_uint159_t(x : std_logic_vector) return uint159_t;
subtype int159_t is signed(158 downto 0);
constant int159_t_SLV_LEN : integer := 159;
function int159_t_to_slv(x : int159_t) return std_logic_vector;
function slv_to_int159_t(x : std_logic_vector) return int159_t;
subtype uint160_t is unsigned(159 downto 0);
constant uint160_t_SLV_LEN : integer := 160;
function uint160_t_to_slv(x : uint160_t) return std_logic_vector;
function slv_to_uint160_t(x : std_logic_vector) return uint160_t;
subtype int160_t is signed(159 downto 0);
constant int160_t_SLV_LEN : integer := 160;
function int160_t_to_slv(x : int160_t) return std_logic_vector;
function slv_to_int160_t(x : std_logic_vector) return int160_t;
subtype uint161_t is unsigned(160 downto 0);
constant uint161_t_SLV_LEN : integer := 161;
function uint161_t_to_slv(x : uint161_t) return std_logic_vector;
function slv_to_uint161_t(x : std_logic_vector) return uint161_t;
subtype int161_t is signed(160 downto 0);
constant int161_t_SLV_LEN : integer := 161;
function int161_t_to_slv(x : int161_t) return std_logic_vector;
function slv_to_int161_t(x : std_logic_vector) return int161_t;
subtype uint162_t is unsigned(161 downto 0);
constant uint162_t_SLV_LEN : integer := 162;
function uint162_t_to_slv(x : uint162_t) return std_logic_vector;
function slv_to_uint162_t(x : std_logic_vector) return uint162_t;
subtype int162_t is signed(161 downto 0);
constant int162_t_SLV_LEN : integer := 162;
function int162_t_to_slv(x : int162_t) return std_logic_vector;
function slv_to_int162_t(x : std_logic_vector) return int162_t;
subtype uint163_t is unsigned(162 downto 0);
constant uint163_t_SLV_LEN : integer := 163;
function uint163_t_to_slv(x : uint163_t) return std_logic_vector;
function slv_to_uint163_t(x : std_logic_vector) return uint163_t;
subtype int163_t is signed(162 downto 0);
constant int163_t_SLV_LEN : integer := 163;
function int163_t_to_slv(x : int163_t) return std_logic_vector;
function slv_to_int163_t(x : std_logic_vector) return int163_t;
subtype uint164_t is unsigned(163 downto 0);
constant uint164_t_SLV_LEN : integer := 164;
function uint164_t_to_slv(x : uint164_t) return std_logic_vector;
function slv_to_uint164_t(x : std_logic_vector) return uint164_t;
subtype int164_t is signed(163 downto 0);
constant int164_t_SLV_LEN : integer := 164;
function int164_t_to_slv(x : int164_t) return std_logic_vector;
function slv_to_int164_t(x : std_logic_vector) return int164_t;
subtype uint165_t is unsigned(164 downto 0);
constant uint165_t_SLV_LEN : integer := 165;
function uint165_t_to_slv(x : uint165_t) return std_logic_vector;
function slv_to_uint165_t(x : std_logic_vector) return uint165_t;
subtype int165_t is signed(164 downto 0);
constant int165_t_SLV_LEN : integer := 165;
function int165_t_to_slv(x : int165_t) return std_logic_vector;
function slv_to_int165_t(x : std_logic_vector) return int165_t;
subtype uint166_t is unsigned(165 downto 0);
constant uint166_t_SLV_LEN : integer := 166;
function uint166_t_to_slv(x : uint166_t) return std_logic_vector;
function slv_to_uint166_t(x : std_logic_vector) return uint166_t;
subtype int166_t is signed(165 downto 0);
constant int166_t_SLV_LEN : integer := 166;
function int166_t_to_slv(x : int166_t) return std_logic_vector;
function slv_to_int166_t(x : std_logic_vector) return int166_t;
subtype uint167_t is unsigned(166 downto 0);
constant uint167_t_SLV_LEN : integer := 167;
function uint167_t_to_slv(x : uint167_t) return std_logic_vector;
function slv_to_uint167_t(x : std_logic_vector) return uint167_t;
subtype int167_t is signed(166 downto 0);
constant int167_t_SLV_LEN : integer := 167;
function int167_t_to_slv(x : int167_t) return std_logic_vector;
function slv_to_int167_t(x : std_logic_vector) return int167_t;
subtype uint168_t is unsigned(167 downto 0);
constant uint168_t_SLV_LEN : integer := 168;
function uint168_t_to_slv(x : uint168_t) return std_logic_vector;
function slv_to_uint168_t(x : std_logic_vector) return uint168_t;
subtype int168_t is signed(167 downto 0);
constant int168_t_SLV_LEN : integer := 168;
function int168_t_to_slv(x : int168_t) return std_logic_vector;
function slv_to_int168_t(x : std_logic_vector) return int168_t;
subtype uint169_t is unsigned(168 downto 0);
constant uint169_t_SLV_LEN : integer := 169;
function uint169_t_to_slv(x : uint169_t) return std_logic_vector;
function slv_to_uint169_t(x : std_logic_vector) return uint169_t;
subtype int169_t is signed(168 downto 0);
constant int169_t_SLV_LEN : integer := 169;
function int169_t_to_slv(x : int169_t) return std_logic_vector;
function slv_to_int169_t(x : std_logic_vector) return int169_t;
subtype uint170_t is unsigned(169 downto 0);
constant uint170_t_SLV_LEN : integer := 170;
function uint170_t_to_slv(x : uint170_t) return std_logic_vector;
function slv_to_uint170_t(x : std_logic_vector) return uint170_t;
subtype int170_t is signed(169 downto 0);
constant int170_t_SLV_LEN : integer := 170;
function int170_t_to_slv(x : int170_t) return std_logic_vector;
function slv_to_int170_t(x : std_logic_vector) return int170_t;
subtype uint171_t is unsigned(170 downto 0);
constant uint171_t_SLV_LEN : integer := 171;
function uint171_t_to_slv(x : uint171_t) return std_logic_vector;
function slv_to_uint171_t(x : std_logic_vector) return uint171_t;
subtype int171_t is signed(170 downto 0);
constant int171_t_SLV_LEN : integer := 171;
function int171_t_to_slv(x : int171_t) return std_logic_vector;
function slv_to_int171_t(x : std_logic_vector) return int171_t;
subtype uint172_t is unsigned(171 downto 0);
constant uint172_t_SLV_LEN : integer := 172;
function uint172_t_to_slv(x : uint172_t) return std_logic_vector;
function slv_to_uint172_t(x : std_logic_vector) return uint172_t;
subtype int172_t is signed(171 downto 0);
constant int172_t_SLV_LEN : integer := 172;
function int172_t_to_slv(x : int172_t) return std_logic_vector;
function slv_to_int172_t(x : std_logic_vector) return int172_t;
subtype uint173_t is unsigned(172 downto 0);
constant uint173_t_SLV_LEN : integer := 173;
function uint173_t_to_slv(x : uint173_t) return std_logic_vector;
function slv_to_uint173_t(x : std_logic_vector) return uint173_t;
subtype int173_t is signed(172 downto 0);
constant int173_t_SLV_LEN : integer := 173;
function int173_t_to_slv(x : int173_t) return std_logic_vector;
function slv_to_int173_t(x : std_logic_vector) return int173_t;
subtype uint174_t is unsigned(173 downto 0);
constant uint174_t_SLV_LEN : integer := 174;
function uint174_t_to_slv(x : uint174_t) return std_logic_vector;
function slv_to_uint174_t(x : std_logic_vector) return uint174_t;
subtype int174_t is signed(173 downto 0);
constant int174_t_SLV_LEN : integer := 174;
function int174_t_to_slv(x : int174_t) return std_logic_vector;
function slv_to_int174_t(x : std_logic_vector) return int174_t;
subtype uint175_t is unsigned(174 downto 0);
constant uint175_t_SLV_LEN : integer := 175;
function uint175_t_to_slv(x : uint175_t) return std_logic_vector;
function slv_to_uint175_t(x : std_logic_vector) return uint175_t;
subtype int175_t is signed(174 downto 0);
constant int175_t_SLV_LEN : integer := 175;
function int175_t_to_slv(x : int175_t) return std_logic_vector;
function slv_to_int175_t(x : std_logic_vector) return int175_t;
subtype uint176_t is unsigned(175 downto 0);
constant uint176_t_SLV_LEN : integer := 176;
function uint176_t_to_slv(x : uint176_t) return std_logic_vector;
function slv_to_uint176_t(x : std_logic_vector) return uint176_t;
subtype int176_t is signed(175 downto 0);
constant int176_t_SLV_LEN : integer := 176;
function int176_t_to_slv(x : int176_t) return std_logic_vector;
function slv_to_int176_t(x : std_logic_vector) return int176_t;
subtype uint177_t is unsigned(176 downto 0);
constant uint177_t_SLV_LEN : integer := 177;
function uint177_t_to_slv(x : uint177_t) return std_logic_vector;
function slv_to_uint177_t(x : std_logic_vector) return uint177_t;
subtype int177_t is signed(176 downto 0);
constant int177_t_SLV_LEN : integer := 177;
function int177_t_to_slv(x : int177_t) return std_logic_vector;
function slv_to_int177_t(x : std_logic_vector) return int177_t;
subtype uint178_t is unsigned(177 downto 0);
constant uint178_t_SLV_LEN : integer := 178;
function uint178_t_to_slv(x : uint178_t) return std_logic_vector;
function slv_to_uint178_t(x : std_logic_vector) return uint178_t;
subtype int178_t is signed(177 downto 0);
constant int178_t_SLV_LEN : integer := 178;
function int178_t_to_slv(x : int178_t) return std_logic_vector;
function slv_to_int178_t(x : std_logic_vector) return int178_t;
subtype uint179_t is unsigned(178 downto 0);
constant uint179_t_SLV_LEN : integer := 179;
function uint179_t_to_slv(x : uint179_t) return std_logic_vector;
function slv_to_uint179_t(x : std_logic_vector) return uint179_t;
subtype int179_t is signed(178 downto 0);
constant int179_t_SLV_LEN : integer := 179;
function int179_t_to_slv(x : int179_t) return std_logic_vector;
function slv_to_int179_t(x : std_logic_vector) return int179_t;
subtype uint180_t is unsigned(179 downto 0);
constant uint180_t_SLV_LEN : integer := 180;
function uint180_t_to_slv(x : uint180_t) return std_logic_vector;
function slv_to_uint180_t(x : std_logic_vector) return uint180_t;
subtype int180_t is signed(179 downto 0);
constant int180_t_SLV_LEN : integer := 180;
function int180_t_to_slv(x : int180_t) return std_logic_vector;
function slv_to_int180_t(x : std_logic_vector) return int180_t;
subtype uint181_t is unsigned(180 downto 0);
constant uint181_t_SLV_LEN : integer := 181;
function uint181_t_to_slv(x : uint181_t) return std_logic_vector;
function slv_to_uint181_t(x : std_logic_vector) return uint181_t;
subtype int181_t is signed(180 downto 0);
constant int181_t_SLV_LEN : integer := 181;
function int181_t_to_slv(x : int181_t) return std_logic_vector;
function slv_to_int181_t(x : std_logic_vector) return int181_t;
subtype uint182_t is unsigned(181 downto 0);
constant uint182_t_SLV_LEN : integer := 182;
function uint182_t_to_slv(x : uint182_t) return std_logic_vector;
function slv_to_uint182_t(x : std_logic_vector) return uint182_t;
subtype int182_t is signed(181 downto 0);
constant int182_t_SLV_LEN : integer := 182;
function int182_t_to_slv(x : int182_t) return std_logic_vector;
function slv_to_int182_t(x : std_logic_vector) return int182_t;
subtype uint183_t is unsigned(182 downto 0);
constant uint183_t_SLV_LEN : integer := 183;
function uint183_t_to_slv(x : uint183_t) return std_logic_vector;
function slv_to_uint183_t(x : std_logic_vector) return uint183_t;
subtype int183_t is signed(182 downto 0);
constant int183_t_SLV_LEN : integer := 183;
function int183_t_to_slv(x : int183_t) return std_logic_vector;
function slv_to_int183_t(x : std_logic_vector) return int183_t;
subtype uint184_t is unsigned(183 downto 0);
constant uint184_t_SLV_LEN : integer := 184;
function uint184_t_to_slv(x : uint184_t) return std_logic_vector;
function slv_to_uint184_t(x : std_logic_vector) return uint184_t;
subtype int184_t is signed(183 downto 0);
constant int184_t_SLV_LEN : integer := 184;
function int184_t_to_slv(x : int184_t) return std_logic_vector;
function slv_to_int184_t(x : std_logic_vector) return int184_t;
subtype uint185_t is unsigned(184 downto 0);
constant uint185_t_SLV_LEN : integer := 185;
function uint185_t_to_slv(x : uint185_t) return std_logic_vector;
function slv_to_uint185_t(x : std_logic_vector) return uint185_t;
subtype int185_t is signed(184 downto 0);
constant int185_t_SLV_LEN : integer := 185;
function int185_t_to_slv(x : int185_t) return std_logic_vector;
function slv_to_int185_t(x : std_logic_vector) return int185_t;
subtype uint186_t is unsigned(185 downto 0);
constant uint186_t_SLV_LEN : integer := 186;
function uint186_t_to_slv(x : uint186_t) return std_logic_vector;
function slv_to_uint186_t(x : std_logic_vector) return uint186_t;
subtype int186_t is signed(185 downto 0);
constant int186_t_SLV_LEN : integer := 186;
function int186_t_to_slv(x : int186_t) return std_logic_vector;
function slv_to_int186_t(x : std_logic_vector) return int186_t;
subtype uint187_t is unsigned(186 downto 0);
constant uint187_t_SLV_LEN : integer := 187;
function uint187_t_to_slv(x : uint187_t) return std_logic_vector;
function slv_to_uint187_t(x : std_logic_vector) return uint187_t;
subtype int187_t is signed(186 downto 0);
constant int187_t_SLV_LEN : integer := 187;
function int187_t_to_slv(x : int187_t) return std_logic_vector;
function slv_to_int187_t(x : std_logic_vector) return int187_t;
subtype uint188_t is unsigned(187 downto 0);
constant uint188_t_SLV_LEN : integer := 188;
function uint188_t_to_slv(x : uint188_t) return std_logic_vector;
function slv_to_uint188_t(x : std_logic_vector) return uint188_t;
subtype int188_t is signed(187 downto 0);
constant int188_t_SLV_LEN : integer := 188;
function int188_t_to_slv(x : int188_t) return std_logic_vector;
function slv_to_int188_t(x : std_logic_vector) return int188_t;
subtype uint189_t is unsigned(188 downto 0);
constant uint189_t_SLV_LEN : integer := 189;
function uint189_t_to_slv(x : uint189_t) return std_logic_vector;
function slv_to_uint189_t(x : std_logic_vector) return uint189_t;
subtype int189_t is signed(188 downto 0);
constant int189_t_SLV_LEN : integer := 189;
function int189_t_to_slv(x : int189_t) return std_logic_vector;
function slv_to_int189_t(x : std_logic_vector) return int189_t;
subtype uint190_t is unsigned(189 downto 0);
constant uint190_t_SLV_LEN : integer := 190;
function uint190_t_to_slv(x : uint190_t) return std_logic_vector;
function slv_to_uint190_t(x : std_logic_vector) return uint190_t;
subtype int190_t is signed(189 downto 0);
constant int190_t_SLV_LEN : integer := 190;
function int190_t_to_slv(x : int190_t) return std_logic_vector;
function slv_to_int190_t(x : std_logic_vector) return int190_t;
subtype uint191_t is unsigned(190 downto 0);
constant uint191_t_SLV_LEN : integer := 191;
function uint191_t_to_slv(x : uint191_t) return std_logic_vector;
function slv_to_uint191_t(x : std_logic_vector) return uint191_t;
subtype int191_t is signed(190 downto 0);
constant int191_t_SLV_LEN : integer := 191;
function int191_t_to_slv(x : int191_t) return std_logic_vector;
function slv_to_int191_t(x : std_logic_vector) return int191_t;
subtype uint192_t is unsigned(191 downto 0);
constant uint192_t_SLV_LEN : integer := 192;
function uint192_t_to_slv(x : uint192_t) return std_logic_vector;
function slv_to_uint192_t(x : std_logic_vector) return uint192_t;
subtype int192_t is signed(191 downto 0);
constant int192_t_SLV_LEN : integer := 192;
function int192_t_to_slv(x : int192_t) return std_logic_vector;
function slv_to_int192_t(x : std_logic_vector) return int192_t;
subtype uint193_t is unsigned(192 downto 0);
constant uint193_t_SLV_LEN : integer := 193;
function uint193_t_to_slv(x : uint193_t) return std_logic_vector;
function slv_to_uint193_t(x : std_logic_vector) return uint193_t;
subtype int193_t is signed(192 downto 0);
constant int193_t_SLV_LEN : integer := 193;
function int193_t_to_slv(x : int193_t) return std_logic_vector;
function slv_to_int193_t(x : std_logic_vector) return int193_t;
subtype uint194_t is unsigned(193 downto 0);
constant uint194_t_SLV_LEN : integer := 194;
function uint194_t_to_slv(x : uint194_t) return std_logic_vector;
function slv_to_uint194_t(x : std_logic_vector) return uint194_t;
subtype int194_t is signed(193 downto 0);
constant int194_t_SLV_LEN : integer := 194;
function int194_t_to_slv(x : int194_t) return std_logic_vector;
function slv_to_int194_t(x : std_logic_vector) return int194_t;
subtype uint195_t is unsigned(194 downto 0);
constant uint195_t_SLV_LEN : integer := 195;
function uint195_t_to_slv(x : uint195_t) return std_logic_vector;
function slv_to_uint195_t(x : std_logic_vector) return uint195_t;
subtype int195_t is signed(194 downto 0);
constant int195_t_SLV_LEN : integer := 195;
function int195_t_to_slv(x : int195_t) return std_logic_vector;
function slv_to_int195_t(x : std_logic_vector) return int195_t;
subtype uint196_t is unsigned(195 downto 0);
constant uint196_t_SLV_LEN : integer := 196;
function uint196_t_to_slv(x : uint196_t) return std_logic_vector;
function slv_to_uint196_t(x : std_logic_vector) return uint196_t;
subtype int196_t is signed(195 downto 0);
constant int196_t_SLV_LEN : integer := 196;
function int196_t_to_slv(x : int196_t) return std_logic_vector;
function slv_to_int196_t(x : std_logic_vector) return int196_t;
subtype uint197_t is unsigned(196 downto 0);
constant uint197_t_SLV_LEN : integer := 197;
function uint197_t_to_slv(x : uint197_t) return std_logic_vector;
function slv_to_uint197_t(x : std_logic_vector) return uint197_t;
subtype int197_t is signed(196 downto 0);
constant int197_t_SLV_LEN : integer := 197;
function int197_t_to_slv(x : int197_t) return std_logic_vector;
function slv_to_int197_t(x : std_logic_vector) return int197_t;
subtype uint198_t is unsigned(197 downto 0);
constant uint198_t_SLV_LEN : integer := 198;
function uint198_t_to_slv(x : uint198_t) return std_logic_vector;
function slv_to_uint198_t(x : std_logic_vector) return uint198_t;
subtype int198_t is signed(197 downto 0);
constant int198_t_SLV_LEN : integer := 198;
function int198_t_to_slv(x : int198_t) return std_logic_vector;
function slv_to_int198_t(x : std_logic_vector) return int198_t;
subtype uint199_t is unsigned(198 downto 0);
constant uint199_t_SLV_LEN : integer := 199;
function uint199_t_to_slv(x : uint199_t) return std_logic_vector;
function slv_to_uint199_t(x : std_logic_vector) return uint199_t;
subtype int199_t is signed(198 downto 0);
constant int199_t_SLV_LEN : integer := 199;
function int199_t_to_slv(x : int199_t) return std_logic_vector;
function slv_to_int199_t(x : std_logic_vector) return int199_t;
subtype uint200_t is unsigned(199 downto 0);
constant uint200_t_SLV_LEN : integer := 200;
function uint200_t_to_slv(x : uint200_t) return std_logic_vector;
function slv_to_uint200_t(x : std_logic_vector) return uint200_t;
subtype int200_t is signed(199 downto 0);
constant int200_t_SLV_LEN : integer := 200;
function int200_t_to_slv(x : int200_t) return std_logic_vector;
function slv_to_int200_t(x : std_logic_vector) return int200_t;
subtype uint201_t is unsigned(200 downto 0);
constant uint201_t_SLV_LEN : integer := 201;
function uint201_t_to_slv(x : uint201_t) return std_logic_vector;
function slv_to_uint201_t(x : std_logic_vector) return uint201_t;
subtype int201_t is signed(200 downto 0);
constant int201_t_SLV_LEN : integer := 201;
function int201_t_to_slv(x : int201_t) return std_logic_vector;
function slv_to_int201_t(x : std_logic_vector) return int201_t;
subtype uint202_t is unsigned(201 downto 0);
constant uint202_t_SLV_LEN : integer := 202;
function uint202_t_to_slv(x : uint202_t) return std_logic_vector;
function slv_to_uint202_t(x : std_logic_vector) return uint202_t;
subtype int202_t is signed(201 downto 0);
constant int202_t_SLV_LEN : integer := 202;
function int202_t_to_slv(x : int202_t) return std_logic_vector;
function slv_to_int202_t(x : std_logic_vector) return int202_t;
subtype uint203_t is unsigned(202 downto 0);
constant uint203_t_SLV_LEN : integer := 203;
function uint203_t_to_slv(x : uint203_t) return std_logic_vector;
function slv_to_uint203_t(x : std_logic_vector) return uint203_t;
subtype int203_t is signed(202 downto 0);
constant int203_t_SLV_LEN : integer := 203;
function int203_t_to_slv(x : int203_t) return std_logic_vector;
function slv_to_int203_t(x : std_logic_vector) return int203_t;
subtype uint204_t is unsigned(203 downto 0);
constant uint204_t_SLV_LEN : integer := 204;
function uint204_t_to_slv(x : uint204_t) return std_logic_vector;
function slv_to_uint204_t(x : std_logic_vector) return uint204_t;
subtype int204_t is signed(203 downto 0);
constant int204_t_SLV_LEN : integer := 204;
function int204_t_to_slv(x : int204_t) return std_logic_vector;
function slv_to_int204_t(x : std_logic_vector) return int204_t;
subtype uint205_t is unsigned(204 downto 0);
constant uint205_t_SLV_LEN : integer := 205;
function uint205_t_to_slv(x : uint205_t) return std_logic_vector;
function slv_to_uint205_t(x : std_logic_vector) return uint205_t;
subtype int205_t is signed(204 downto 0);
constant int205_t_SLV_LEN : integer := 205;
function int205_t_to_slv(x : int205_t) return std_logic_vector;
function slv_to_int205_t(x : std_logic_vector) return int205_t;
subtype uint206_t is unsigned(205 downto 0);
constant uint206_t_SLV_LEN : integer := 206;
function uint206_t_to_slv(x : uint206_t) return std_logic_vector;
function slv_to_uint206_t(x : std_logic_vector) return uint206_t;
subtype int206_t is signed(205 downto 0);
constant int206_t_SLV_LEN : integer := 206;
function int206_t_to_slv(x : int206_t) return std_logic_vector;
function slv_to_int206_t(x : std_logic_vector) return int206_t;
subtype uint207_t is unsigned(206 downto 0);
constant uint207_t_SLV_LEN : integer := 207;
function uint207_t_to_slv(x : uint207_t) return std_logic_vector;
function slv_to_uint207_t(x : std_logic_vector) return uint207_t;
subtype int207_t is signed(206 downto 0);
constant int207_t_SLV_LEN : integer := 207;
function int207_t_to_slv(x : int207_t) return std_logic_vector;
function slv_to_int207_t(x : std_logic_vector) return int207_t;
subtype uint208_t is unsigned(207 downto 0);
constant uint208_t_SLV_LEN : integer := 208;
function uint208_t_to_slv(x : uint208_t) return std_logic_vector;
function slv_to_uint208_t(x : std_logic_vector) return uint208_t;
subtype int208_t is signed(207 downto 0);
constant int208_t_SLV_LEN : integer := 208;
function int208_t_to_slv(x : int208_t) return std_logic_vector;
function slv_to_int208_t(x : std_logic_vector) return int208_t;
subtype uint209_t is unsigned(208 downto 0);
constant uint209_t_SLV_LEN : integer := 209;
function uint209_t_to_slv(x : uint209_t) return std_logic_vector;
function slv_to_uint209_t(x : std_logic_vector) return uint209_t;
subtype int209_t is signed(208 downto 0);
constant int209_t_SLV_LEN : integer := 209;
function int209_t_to_slv(x : int209_t) return std_logic_vector;
function slv_to_int209_t(x : std_logic_vector) return int209_t;
subtype uint210_t is unsigned(209 downto 0);
constant uint210_t_SLV_LEN : integer := 210;
function uint210_t_to_slv(x : uint210_t) return std_logic_vector;
function slv_to_uint210_t(x : std_logic_vector) return uint210_t;
subtype int210_t is signed(209 downto 0);
constant int210_t_SLV_LEN : integer := 210;
function int210_t_to_slv(x : int210_t) return std_logic_vector;
function slv_to_int210_t(x : std_logic_vector) return int210_t;
subtype uint211_t is unsigned(210 downto 0);
constant uint211_t_SLV_LEN : integer := 211;
function uint211_t_to_slv(x : uint211_t) return std_logic_vector;
function slv_to_uint211_t(x : std_logic_vector) return uint211_t;
subtype int211_t is signed(210 downto 0);
constant int211_t_SLV_LEN : integer := 211;
function int211_t_to_slv(x : int211_t) return std_logic_vector;
function slv_to_int211_t(x : std_logic_vector) return int211_t;
subtype uint212_t is unsigned(211 downto 0);
constant uint212_t_SLV_LEN : integer := 212;
function uint212_t_to_slv(x : uint212_t) return std_logic_vector;
function slv_to_uint212_t(x : std_logic_vector) return uint212_t;
subtype int212_t is signed(211 downto 0);
constant int212_t_SLV_LEN : integer := 212;
function int212_t_to_slv(x : int212_t) return std_logic_vector;
function slv_to_int212_t(x : std_logic_vector) return int212_t;
subtype uint213_t is unsigned(212 downto 0);
constant uint213_t_SLV_LEN : integer := 213;
function uint213_t_to_slv(x : uint213_t) return std_logic_vector;
function slv_to_uint213_t(x : std_logic_vector) return uint213_t;
subtype int213_t is signed(212 downto 0);
constant int213_t_SLV_LEN : integer := 213;
function int213_t_to_slv(x : int213_t) return std_logic_vector;
function slv_to_int213_t(x : std_logic_vector) return int213_t;
subtype uint214_t is unsigned(213 downto 0);
constant uint214_t_SLV_LEN : integer := 214;
function uint214_t_to_slv(x : uint214_t) return std_logic_vector;
function slv_to_uint214_t(x : std_logic_vector) return uint214_t;
subtype int214_t is signed(213 downto 0);
constant int214_t_SLV_LEN : integer := 214;
function int214_t_to_slv(x : int214_t) return std_logic_vector;
function slv_to_int214_t(x : std_logic_vector) return int214_t;
subtype uint215_t is unsigned(214 downto 0);
constant uint215_t_SLV_LEN : integer := 215;
function uint215_t_to_slv(x : uint215_t) return std_logic_vector;
function slv_to_uint215_t(x : std_logic_vector) return uint215_t;
subtype int215_t is signed(214 downto 0);
constant int215_t_SLV_LEN : integer := 215;
function int215_t_to_slv(x : int215_t) return std_logic_vector;
function slv_to_int215_t(x : std_logic_vector) return int215_t;
subtype uint216_t is unsigned(215 downto 0);
constant uint216_t_SLV_LEN : integer := 216;
function uint216_t_to_slv(x : uint216_t) return std_logic_vector;
function slv_to_uint216_t(x : std_logic_vector) return uint216_t;
subtype int216_t is signed(215 downto 0);
constant int216_t_SLV_LEN : integer := 216;
function int216_t_to_slv(x : int216_t) return std_logic_vector;
function slv_to_int216_t(x : std_logic_vector) return int216_t;
subtype uint217_t is unsigned(216 downto 0);
constant uint217_t_SLV_LEN : integer := 217;
function uint217_t_to_slv(x : uint217_t) return std_logic_vector;
function slv_to_uint217_t(x : std_logic_vector) return uint217_t;
subtype int217_t is signed(216 downto 0);
constant int217_t_SLV_LEN : integer := 217;
function int217_t_to_slv(x : int217_t) return std_logic_vector;
function slv_to_int217_t(x : std_logic_vector) return int217_t;
subtype uint218_t is unsigned(217 downto 0);
constant uint218_t_SLV_LEN : integer := 218;
function uint218_t_to_slv(x : uint218_t) return std_logic_vector;
function slv_to_uint218_t(x : std_logic_vector) return uint218_t;
subtype int218_t is signed(217 downto 0);
constant int218_t_SLV_LEN : integer := 218;
function int218_t_to_slv(x : int218_t) return std_logic_vector;
function slv_to_int218_t(x : std_logic_vector) return int218_t;
subtype uint219_t is unsigned(218 downto 0);
constant uint219_t_SLV_LEN : integer := 219;
function uint219_t_to_slv(x : uint219_t) return std_logic_vector;
function slv_to_uint219_t(x : std_logic_vector) return uint219_t;
subtype int219_t is signed(218 downto 0);
constant int219_t_SLV_LEN : integer := 219;
function int219_t_to_slv(x : int219_t) return std_logic_vector;
function slv_to_int219_t(x : std_logic_vector) return int219_t;
subtype uint220_t is unsigned(219 downto 0);
constant uint220_t_SLV_LEN : integer := 220;
function uint220_t_to_slv(x : uint220_t) return std_logic_vector;
function slv_to_uint220_t(x : std_logic_vector) return uint220_t;
subtype int220_t is signed(219 downto 0);
constant int220_t_SLV_LEN : integer := 220;
function int220_t_to_slv(x : int220_t) return std_logic_vector;
function slv_to_int220_t(x : std_logic_vector) return int220_t;
subtype uint221_t is unsigned(220 downto 0);
constant uint221_t_SLV_LEN : integer := 221;
function uint221_t_to_slv(x : uint221_t) return std_logic_vector;
function slv_to_uint221_t(x : std_logic_vector) return uint221_t;
subtype int221_t is signed(220 downto 0);
constant int221_t_SLV_LEN : integer := 221;
function int221_t_to_slv(x : int221_t) return std_logic_vector;
function slv_to_int221_t(x : std_logic_vector) return int221_t;
subtype uint222_t is unsigned(221 downto 0);
constant uint222_t_SLV_LEN : integer := 222;
function uint222_t_to_slv(x : uint222_t) return std_logic_vector;
function slv_to_uint222_t(x : std_logic_vector) return uint222_t;
subtype int222_t is signed(221 downto 0);
constant int222_t_SLV_LEN : integer := 222;
function int222_t_to_slv(x : int222_t) return std_logic_vector;
function slv_to_int222_t(x : std_logic_vector) return int222_t;
subtype uint223_t is unsigned(222 downto 0);
constant uint223_t_SLV_LEN : integer := 223;
function uint223_t_to_slv(x : uint223_t) return std_logic_vector;
function slv_to_uint223_t(x : std_logic_vector) return uint223_t;
subtype int223_t is signed(222 downto 0);
constant int223_t_SLV_LEN : integer := 223;
function int223_t_to_slv(x : int223_t) return std_logic_vector;
function slv_to_int223_t(x : std_logic_vector) return int223_t;
subtype uint224_t is unsigned(223 downto 0);
constant uint224_t_SLV_LEN : integer := 224;
function uint224_t_to_slv(x : uint224_t) return std_logic_vector;
function slv_to_uint224_t(x : std_logic_vector) return uint224_t;
subtype int224_t is signed(223 downto 0);
constant int224_t_SLV_LEN : integer := 224;
function int224_t_to_slv(x : int224_t) return std_logic_vector;
function slv_to_int224_t(x : std_logic_vector) return int224_t;
subtype uint225_t is unsigned(224 downto 0);
constant uint225_t_SLV_LEN : integer := 225;
function uint225_t_to_slv(x : uint225_t) return std_logic_vector;
function slv_to_uint225_t(x : std_logic_vector) return uint225_t;
subtype int225_t is signed(224 downto 0);
constant int225_t_SLV_LEN : integer := 225;
function int225_t_to_slv(x : int225_t) return std_logic_vector;
function slv_to_int225_t(x : std_logic_vector) return int225_t;
subtype uint226_t is unsigned(225 downto 0);
constant uint226_t_SLV_LEN : integer := 226;
function uint226_t_to_slv(x : uint226_t) return std_logic_vector;
function slv_to_uint226_t(x : std_logic_vector) return uint226_t;
subtype int226_t is signed(225 downto 0);
constant int226_t_SLV_LEN : integer := 226;
function int226_t_to_slv(x : int226_t) return std_logic_vector;
function slv_to_int226_t(x : std_logic_vector) return int226_t;
subtype uint227_t is unsigned(226 downto 0);
constant uint227_t_SLV_LEN : integer := 227;
function uint227_t_to_slv(x : uint227_t) return std_logic_vector;
function slv_to_uint227_t(x : std_logic_vector) return uint227_t;
subtype int227_t is signed(226 downto 0);
constant int227_t_SLV_LEN : integer := 227;
function int227_t_to_slv(x : int227_t) return std_logic_vector;
function slv_to_int227_t(x : std_logic_vector) return int227_t;
subtype uint228_t is unsigned(227 downto 0);
constant uint228_t_SLV_LEN : integer := 228;
function uint228_t_to_slv(x : uint228_t) return std_logic_vector;
function slv_to_uint228_t(x : std_logic_vector) return uint228_t;
subtype int228_t is signed(227 downto 0);
constant int228_t_SLV_LEN : integer := 228;
function int228_t_to_slv(x : int228_t) return std_logic_vector;
function slv_to_int228_t(x : std_logic_vector) return int228_t;
subtype uint229_t is unsigned(228 downto 0);
constant uint229_t_SLV_LEN : integer := 229;
function uint229_t_to_slv(x : uint229_t) return std_logic_vector;
function slv_to_uint229_t(x : std_logic_vector) return uint229_t;
subtype int229_t is signed(228 downto 0);
constant int229_t_SLV_LEN : integer := 229;
function int229_t_to_slv(x : int229_t) return std_logic_vector;
function slv_to_int229_t(x : std_logic_vector) return int229_t;
subtype uint230_t is unsigned(229 downto 0);
constant uint230_t_SLV_LEN : integer := 230;
function uint230_t_to_slv(x : uint230_t) return std_logic_vector;
function slv_to_uint230_t(x : std_logic_vector) return uint230_t;
subtype int230_t is signed(229 downto 0);
constant int230_t_SLV_LEN : integer := 230;
function int230_t_to_slv(x : int230_t) return std_logic_vector;
function slv_to_int230_t(x : std_logic_vector) return int230_t;
subtype uint231_t is unsigned(230 downto 0);
constant uint231_t_SLV_LEN : integer := 231;
function uint231_t_to_slv(x : uint231_t) return std_logic_vector;
function slv_to_uint231_t(x : std_logic_vector) return uint231_t;
subtype int231_t is signed(230 downto 0);
constant int231_t_SLV_LEN : integer := 231;
function int231_t_to_slv(x : int231_t) return std_logic_vector;
function slv_to_int231_t(x : std_logic_vector) return int231_t;
subtype uint232_t is unsigned(231 downto 0);
constant uint232_t_SLV_LEN : integer := 232;
function uint232_t_to_slv(x : uint232_t) return std_logic_vector;
function slv_to_uint232_t(x : std_logic_vector) return uint232_t;
subtype int232_t is signed(231 downto 0);
constant int232_t_SLV_LEN : integer := 232;
function int232_t_to_slv(x : int232_t) return std_logic_vector;
function slv_to_int232_t(x : std_logic_vector) return int232_t;
subtype uint233_t is unsigned(232 downto 0);
constant uint233_t_SLV_LEN : integer := 233;
function uint233_t_to_slv(x : uint233_t) return std_logic_vector;
function slv_to_uint233_t(x : std_logic_vector) return uint233_t;
subtype int233_t is signed(232 downto 0);
constant int233_t_SLV_LEN : integer := 233;
function int233_t_to_slv(x : int233_t) return std_logic_vector;
function slv_to_int233_t(x : std_logic_vector) return int233_t;
subtype uint234_t is unsigned(233 downto 0);
constant uint234_t_SLV_LEN : integer := 234;
function uint234_t_to_slv(x : uint234_t) return std_logic_vector;
function slv_to_uint234_t(x : std_logic_vector) return uint234_t;
subtype int234_t is signed(233 downto 0);
constant int234_t_SLV_LEN : integer := 234;
function int234_t_to_slv(x : int234_t) return std_logic_vector;
function slv_to_int234_t(x : std_logic_vector) return int234_t;
subtype uint235_t is unsigned(234 downto 0);
constant uint235_t_SLV_LEN : integer := 235;
function uint235_t_to_slv(x : uint235_t) return std_logic_vector;
function slv_to_uint235_t(x : std_logic_vector) return uint235_t;
subtype int235_t is signed(234 downto 0);
constant int235_t_SLV_LEN : integer := 235;
function int235_t_to_slv(x : int235_t) return std_logic_vector;
function slv_to_int235_t(x : std_logic_vector) return int235_t;
subtype uint236_t is unsigned(235 downto 0);
constant uint236_t_SLV_LEN : integer := 236;
function uint236_t_to_slv(x : uint236_t) return std_logic_vector;
function slv_to_uint236_t(x : std_logic_vector) return uint236_t;
subtype int236_t is signed(235 downto 0);
constant int236_t_SLV_LEN : integer := 236;
function int236_t_to_slv(x : int236_t) return std_logic_vector;
function slv_to_int236_t(x : std_logic_vector) return int236_t;
subtype uint237_t is unsigned(236 downto 0);
constant uint237_t_SLV_LEN : integer := 237;
function uint237_t_to_slv(x : uint237_t) return std_logic_vector;
function slv_to_uint237_t(x : std_logic_vector) return uint237_t;
subtype int237_t is signed(236 downto 0);
constant int237_t_SLV_LEN : integer := 237;
function int237_t_to_slv(x : int237_t) return std_logic_vector;
function slv_to_int237_t(x : std_logic_vector) return int237_t;
subtype uint238_t is unsigned(237 downto 0);
constant uint238_t_SLV_LEN : integer := 238;
function uint238_t_to_slv(x : uint238_t) return std_logic_vector;
function slv_to_uint238_t(x : std_logic_vector) return uint238_t;
subtype int238_t is signed(237 downto 0);
constant int238_t_SLV_LEN : integer := 238;
function int238_t_to_slv(x : int238_t) return std_logic_vector;
function slv_to_int238_t(x : std_logic_vector) return int238_t;
subtype uint239_t is unsigned(238 downto 0);
constant uint239_t_SLV_LEN : integer := 239;
function uint239_t_to_slv(x : uint239_t) return std_logic_vector;
function slv_to_uint239_t(x : std_logic_vector) return uint239_t;
subtype int239_t is signed(238 downto 0);
constant int239_t_SLV_LEN : integer := 239;
function int239_t_to_slv(x : int239_t) return std_logic_vector;
function slv_to_int239_t(x : std_logic_vector) return int239_t;
subtype uint240_t is unsigned(239 downto 0);
constant uint240_t_SLV_LEN : integer := 240;
function uint240_t_to_slv(x : uint240_t) return std_logic_vector;
function slv_to_uint240_t(x : std_logic_vector) return uint240_t;
subtype int240_t is signed(239 downto 0);
constant int240_t_SLV_LEN : integer := 240;
function int240_t_to_slv(x : int240_t) return std_logic_vector;
function slv_to_int240_t(x : std_logic_vector) return int240_t;
subtype uint241_t is unsigned(240 downto 0);
constant uint241_t_SLV_LEN : integer := 241;
function uint241_t_to_slv(x : uint241_t) return std_logic_vector;
function slv_to_uint241_t(x : std_logic_vector) return uint241_t;
subtype int241_t is signed(240 downto 0);
constant int241_t_SLV_LEN : integer := 241;
function int241_t_to_slv(x : int241_t) return std_logic_vector;
function slv_to_int241_t(x : std_logic_vector) return int241_t;
subtype uint242_t is unsigned(241 downto 0);
constant uint242_t_SLV_LEN : integer := 242;
function uint242_t_to_slv(x : uint242_t) return std_logic_vector;
function slv_to_uint242_t(x : std_logic_vector) return uint242_t;
subtype int242_t is signed(241 downto 0);
constant int242_t_SLV_LEN : integer := 242;
function int242_t_to_slv(x : int242_t) return std_logic_vector;
function slv_to_int242_t(x : std_logic_vector) return int242_t;
subtype uint243_t is unsigned(242 downto 0);
constant uint243_t_SLV_LEN : integer := 243;
function uint243_t_to_slv(x : uint243_t) return std_logic_vector;
function slv_to_uint243_t(x : std_logic_vector) return uint243_t;
subtype int243_t is signed(242 downto 0);
constant int243_t_SLV_LEN : integer := 243;
function int243_t_to_slv(x : int243_t) return std_logic_vector;
function slv_to_int243_t(x : std_logic_vector) return int243_t;
subtype uint244_t is unsigned(243 downto 0);
constant uint244_t_SLV_LEN : integer := 244;
function uint244_t_to_slv(x : uint244_t) return std_logic_vector;
function slv_to_uint244_t(x : std_logic_vector) return uint244_t;
subtype int244_t is signed(243 downto 0);
constant int244_t_SLV_LEN : integer := 244;
function int244_t_to_slv(x : int244_t) return std_logic_vector;
function slv_to_int244_t(x : std_logic_vector) return int244_t;
subtype uint245_t is unsigned(244 downto 0);
constant uint245_t_SLV_LEN : integer := 245;
function uint245_t_to_slv(x : uint245_t) return std_logic_vector;
function slv_to_uint245_t(x : std_logic_vector) return uint245_t;
subtype int245_t is signed(244 downto 0);
constant int245_t_SLV_LEN : integer := 245;
function int245_t_to_slv(x : int245_t) return std_logic_vector;
function slv_to_int245_t(x : std_logic_vector) return int245_t;
subtype uint246_t is unsigned(245 downto 0);
constant uint246_t_SLV_LEN : integer := 246;
function uint246_t_to_slv(x : uint246_t) return std_logic_vector;
function slv_to_uint246_t(x : std_logic_vector) return uint246_t;
subtype int246_t is signed(245 downto 0);
constant int246_t_SLV_LEN : integer := 246;
function int246_t_to_slv(x : int246_t) return std_logic_vector;
function slv_to_int246_t(x : std_logic_vector) return int246_t;
subtype uint247_t is unsigned(246 downto 0);
constant uint247_t_SLV_LEN : integer := 247;
function uint247_t_to_slv(x : uint247_t) return std_logic_vector;
function slv_to_uint247_t(x : std_logic_vector) return uint247_t;
subtype int247_t is signed(246 downto 0);
constant int247_t_SLV_LEN : integer := 247;
function int247_t_to_slv(x : int247_t) return std_logic_vector;
function slv_to_int247_t(x : std_logic_vector) return int247_t;
subtype uint248_t is unsigned(247 downto 0);
constant uint248_t_SLV_LEN : integer := 248;
function uint248_t_to_slv(x : uint248_t) return std_logic_vector;
function slv_to_uint248_t(x : std_logic_vector) return uint248_t;
subtype int248_t is signed(247 downto 0);
constant int248_t_SLV_LEN : integer := 248;
function int248_t_to_slv(x : int248_t) return std_logic_vector;
function slv_to_int248_t(x : std_logic_vector) return int248_t;
subtype uint249_t is unsigned(248 downto 0);
constant uint249_t_SLV_LEN : integer := 249;
function uint249_t_to_slv(x : uint249_t) return std_logic_vector;
function slv_to_uint249_t(x : std_logic_vector) return uint249_t;
subtype int249_t is signed(248 downto 0);
constant int249_t_SLV_LEN : integer := 249;
function int249_t_to_slv(x : int249_t) return std_logic_vector;
function slv_to_int249_t(x : std_logic_vector) return int249_t;
subtype uint250_t is unsigned(249 downto 0);
constant uint250_t_SLV_LEN : integer := 250;
function uint250_t_to_slv(x : uint250_t) return std_logic_vector;
function slv_to_uint250_t(x : std_logic_vector) return uint250_t;
subtype int250_t is signed(249 downto 0);
constant int250_t_SLV_LEN : integer := 250;
function int250_t_to_slv(x : int250_t) return std_logic_vector;
function slv_to_int250_t(x : std_logic_vector) return int250_t;
subtype uint251_t is unsigned(250 downto 0);
constant uint251_t_SLV_LEN : integer := 251;
function uint251_t_to_slv(x : uint251_t) return std_logic_vector;
function slv_to_uint251_t(x : std_logic_vector) return uint251_t;
subtype int251_t is signed(250 downto 0);
constant int251_t_SLV_LEN : integer := 251;
function int251_t_to_slv(x : int251_t) return std_logic_vector;
function slv_to_int251_t(x : std_logic_vector) return int251_t;
subtype uint252_t is unsigned(251 downto 0);
constant uint252_t_SLV_LEN : integer := 252;
function uint252_t_to_slv(x : uint252_t) return std_logic_vector;
function slv_to_uint252_t(x : std_logic_vector) return uint252_t;
subtype int252_t is signed(251 downto 0);
constant int252_t_SLV_LEN : integer := 252;
function int252_t_to_slv(x : int252_t) return std_logic_vector;
function slv_to_int252_t(x : std_logic_vector) return int252_t;
subtype uint253_t is unsigned(252 downto 0);
constant uint253_t_SLV_LEN : integer := 253;
function uint253_t_to_slv(x : uint253_t) return std_logic_vector;
function slv_to_uint253_t(x : std_logic_vector) return uint253_t;
subtype int253_t is signed(252 downto 0);
constant int253_t_SLV_LEN : integer := 253;
function int253_t_to_slv(x : int253_t) return std_logic_vector;
function slv_to_int253_t(x : std_logic_vector) return int253_t;
subtype uint254_t is unsigned(253 downto 0);
constant uint254_t_SLV_LEN : integer := 254;
function uint254_t_to_slv(x : uint254_t) return std_logic_vector;
function slv_to_uint254_t(x : std_logic_vector) return uint254_t;
subtype int254_t is signed(253 downto 0);
constant int254_t_SLV_LEN : integer := 254;
function int254_t_to_slv(x : int254_t) return std_logic_vector;
function slv_to_int254_t(x : std_logic_vector) return int254_t;
subtype uint255_t is unsigned(254 downto 0);
constant uint255_t_SLV_LEN : integer := 255;
function uint255_t_to_slv(x : uint255_t) return std_logic_vector;
function slv_to_uint255_t(x : std_logic_vector) return uint255_t;
subtype int255_t is signed(254 downto 0);
constant int255_t_SLV_LEN : integer := 255;
function int255_t_to_slv(x : int255_t) return std_logic_vector;
function slv_to_int255_t(x : std_logic_vector) return int255_t;
subtype uint256_t is unsigned(255 downto 0);
constant uint256_t_SLV_LEN : integer := 256;
function uint256_t_to_slv(x : uint256_t) return std_logic_vector;
function slv_to_uint256_t(x : std_logic_vector) return uint256_t;
subtype int256_t is signed(255 downto 0);
constant int256_t_SLV_LEN : integer := 256;
function int256_t_to_slv(x : int256_t) return std_logic_vector;
function slv_to_int256_t(x : std_logic_vector) return int256_t;
subtype uint257_t is unsigned(256 downto 0);
constant uint257_t_SLV_LEN : integer := 257;
function uint257_t_to_slv(x : uint257_t) return std_logic_vector;
function slv_to_uint257_t(x : std_logic_vector) return uint257_t;
subtype int257_t is signed(256 downto 0);
constant int257_t_SLV_LEN : integer := 257;
function int257_t_to_slv(x : int257_t) return std_logic_vector;
function slv_to_int257_t(x : std_logic_vector) return int257_t;
subtype uint258_t is unsigned(257 downto 0);
constant uint258_t_SLV_LEN : integer := 258;
function uint258_t_to_slv(x : uint258_t) return std_logic_vector;
function slv_to_uint258_t(x : std_logic_vector) return uint258_t;
subtype int258_t is signed(257 downto 0);
constant int258_t_SLV_LEN : integer := 258;
function int258_t_to_slv(x : int258_t) return std_logic_vector;
function slv_to_int258_t(x : std_logic_vector) return int258_t;
subtype uint259_t is unsigned(258 downto 0);
constant uint259_t_SLV_LEN : integer := 259;
function uint259_t_to_slv(x : uint259_t) return std_logic_vector;
function slv_to_uint259_t(x : std_logic_vector) return uint259_t;
subtype int259_t is signed(258 downto 0);
constant int259_t_SLV_LEN : integer := 259;
function int259_t_to_slv(x : int259_t) return std_logic_vector;
function slv_to_int259_t(x : std_logic_vector) return int259_t;
subtype uint260_t is unsigned(259 downto 0);
constant uint260_t_SLV_LEN : integer := 260;
function uint260_t_to_slv(x : uint260_t) return std_logic_vector;
function slv_to_uint260_t(x : std_logic_vector) return uint260_t;
subtype int260_t is signed(259 downto 0);
constant int260_t_SLV_LEN : integer := 260;
function int260_t_to_slv(x : int260_t) return std_logic_vector;
function slv_to_int260_t(x : std_logic_vector) return int260_t;
subtype uint261_t is unsigned(260 downto 0);
constant uint261_t_SLV_LEN : integer := 261;
function uint261_t_to_slv(x : uint261_t) return std_logic_vector;
function slv_to_uint261_t(x : std_logic_vector) return uint261_t;
subtype int261_t is signed(260 downto 0);
constant int261_t_SLV_LEN : integer := 261;
function int261_t_to_slv(x : int261_t) return std_logic_vector;
function slv_to_int261_t(x : std_logic_vector) return int261_t;
subtype uint262_t is unsigned(261 downto 0);
constant uint262_t_SLV_LEN : integer := 262;
function uint262_t_to_slv(x : uint262_t) return std_logic_vector;
function slv_to_uint262_t(x : std_logic_vector) return uint262_t;
subtype int262_t is signed(261 downto 0);
constant int262_t_SLV_LEN : integer := 262;
function int262_t_to_slv(x : int262_t) return std_logic_vector;
function slv_to_int262_t(x : std_logic_vector) return int262_t;
subtype uint263_t is unsigned(262 downto 0);
constant uint263_t_SLV_LEN : integer := 263;
function uint263_t_to_slv(x : uint263_t) return std_logic_vector;
function slv_to_uint263_t(x : std_logic_vector) return uint263_t;
subtype int263_t is signed(262 downto 0);
constant int263_t_SLV_LEN : integer := 263;
function int263_t_to_slv(x : int263_t) return std_logic_vector;
function slv_to_int263_t(x : std_logic_vector) return int263_t;
subtype uint264_t is unsigned(263 downto 0);
constant uint264_t_SLV_LEN : integer := 264;
function uint264_t_to_slv(x : uint264_t) return std_logic_vector;
function slv_to_uint264_t(x : std_logic_vector) return uint264_t;
subtype int264_t is signed(263 downto 0);
constant int264_t_SLV_LEN : integer := 264;
function int264_t_to_slv(x : int264_t) return std_logic_vector;
function slv_to_int264_t(x : std_logic_vector) return int264_t;
subtype uint265_t is unsigned(264 downto 0);
constant uint265_t_SLV_LEN : integer := 265;
function uint265_t_to_slv(x : uint265_t) return std_logic_vector;
function slv_to_uint265_t(x : std_logic_vector) return uint265_t;
subtype int265_t is signed(264 downto 0);
constant int265_t_SLV_LEN : integer := 265;
function int265_t_to_slv(x : int265_t) return std_logic_vector;
function slv_to_int265_t(x : std_logic_vector) return int265_t;
subtype uint266_t is unsigned(265 downto 0);
constant uint266_t_SLV_LEN : integer := 266;
function uint266_t_to_slv(x : uint266_t) return std_logic_vector;
function slv_to_uint266_t(x : std_logic_vector) return uint266_t;
subtype int266_t is signed(265 downto 0);
constant int266_t_SLV_LEN : integer := 266;
function int266_t_to_slv(x : int266_t) return std_logic_vector;
function slv_to_int266_t(x : std_logic_vector) return int266_t;
subtype uint267_t is unsigned(266 downto 0);
constant uint267_t_SLV_LEN : integer := 267;
function uint267_t_to_slv(x : uint267_t) return std_logic_vector;
function slv_to_uint267_t(x : std_logic_vector) return uint267_t;
subtype int267_t is signed(266 downto 0);
constant int267_t_SLV_LEN : integer := 267;
function int267_t_to_slv(x : int267_t) return std_logic_vector;
function slv_to_int267_t(x : std_logic_vector) return int267_t;
subtype uint268_t is unsigned(267 downto 0);
constant uint268_t_SLV_LEN : integer := 268;
function uint268_t_to_slv(x : uint268_t) return std_logic_vector;
function slv_to_uint268_t(x : std_logic_vector) return uint268_t;
subtype int268_t is signed(267 downto 0);
constant int268_t_SLV_LEN : integer := 268;
function int268_t_to_slv(x : int268_t) return std_logic_vector;
function slv_to_int268_t(x : std_logic_vector) return int268_t;
subtype uint269_t is unsigned(268 downto 0);
constant uint269_t_SLV_LEN : integer := 269;
function uint269_t_to_slv(x : uint269_t) return std_logic_vector;
function slv_to_uint269_t(x : std_logic_vector) return uint269_t;
subtype int269_t is signed(268 downto 0);
constant int269_t_SLV_LEN : integer := 269;
function int269_t_to_slv(x : int269_t) return std_logic_vector;
function slv_to_int269_t(x : std_logic_vector) return int269_t;
subtype uint270_t is unsigned(269 downto 0);
constant uint270_t_SLV_LEN : integer := 270;
function uint270_t_to_slv(x : uint270_t) return std_logic_vector;
function slv_to_uint270_t(x : std_logic_vector) return uint270_t;
subtype int270_t is signed(269 downto 0);
constant int270_t_SLV_LEN : integer := 270;
function int270_t_to_slv(x : int270_t) return std_logic_vector;
function slv_to_int270_t(x : std_logic_vector) return int270_t;
subtype uint271_t is unsigned(270 downto 0);
constant uint271_t_SLV_LEN : integer := 271;
function uint271_t_to_slv(x : uint271_t) return std_logic_vector;
function slv_to_uint271_t(x : std_logic_vector) return uint271_t;
subtype int271_t is signed(270 downto 0);
constant int271_t_SLV_LEN : integer := 271;
function int271_t_to_slv(x : int271_t) return std_logic_vector;
function slv_to_int271_t(x : std_logic_vector) return int271_t;
subtype uint272_t is unsigned(271 downto 0);
constant uint272_t_SLV_LEN : integer := 272;
function uint272_t_to_slv(x : uint272_t) return std_logic_vector;
function slv_to_uint272_t(x : std_logic_vector) return uint272_t;
subtype int272_t is signed(271 downto 0);
constant int272_t_SLV_LEN : integer := 272;
function int272_t_to_slv(x : int272_t) return std_logic_vector;
function slv_to_int272_t(x : std_logic_vector) return int272_t;
subtype uint273_t is unsigned(272 downto 0);
constant uint273_t_SLV_LEN : integer := 273;
function uint273_t_to_slv(x : uint273_t) return std_logic_vector;
function slv_to_uint273_t(x : std_logic_vector) return uint273_t;
subtype int273_t is signed(272 downto 0);
constant int273_t_SLV_LEN : integer := 273;
function int273_t_to_slv(x : int273_t) return std_logic_vector;
function slv_to_int273_t(x : std_logic_vector) return int273_t;
subtype uint274_t is unsigned(273 downto 0);
constant uint274_t_SLV_LEN : integer := 274;
function uint274_t_to_slv(x : uint274_t) return std_logic_vector;
function slv_to_uint274_t(x : std_logic_vector) return uint274_t;
subtype int274_t is signed(273 downto 0);
constant int274_t_SLV_LEN : integer := 274;
function int274_t_to_slv(x : int274_t) return std_logic_vector;
function slv_to_int274_t(x : std_logic_vector) return int274_t;
subtype uint275_t is unsigned(274 downto 0);
constant uint275_t_SLV_LEN : integer := 275;
function uint275_t_to_slv(x : uint275_t) return std_logic_vector;
function slv_to_uint275_t(x : std_logic_vector) return uint275_t;
subtype int275_t is signed(274 downto 0);
constant int275_t_SLV_LEN : integer := 275;
function int275_t_to_slv(x : int275_t) return std_logic_vector;
function slv_to_int275_t(x : std_logic_vector) return int275_t;
subtype uint276_t is unsigned(275 downto 0);
constant uint276_t_SLV_LEN : integer := 276;
function uint276_t_to_slv(x : uint276_t) return std_logic_vector;
function slv_to_uint276_t(x : std_logic_vector) return uint276_t;
subtype int276_t is signed(275 downto 0);
constant int276_t_SLV_LEN : integer := 276;
function int276_t_to_slv(x : int276_t) return std_logic_vector;
function slv_to_int276_t(x : std_logic_vector) return int276_t;
subtype uint277_t is unsigned(276 downto 0);
constant uint277_t_SLV_LEN : integer := 277;
function uint277_t_to_slv(x : uint277_t) return std_logic_vector;
function slv_to_uint277_t(x : std_logic_vector) return uint277_t;
subtype int277_t is signed(276 downto 0);
constant int277_t_SLV_LEN : integer := 277;
function int277_t_to_slv(x : int277_t) return std_logic_vector;
function slv_to_int277_t(x : std_logic_vector) return int277_t;
subtype uint278_t is unsigned(277 downto 0);
constant uint278_t_SLV_LEN : integer := 278;
function uint278_t_to_slv(x : uint278_t) return std_logic_vector;
function slv_to_uint278_t(x : std_logic_vector) return uint278_t;
subtype int278_t is signed(277 downto 0);
constant int278_t_SLV_LEN : integer := 278;
function int278_t_to_slv(x : int278_t) return std_logic_vector;
function slv_to_int278_t(x : std_logic_vector) return int278_t;
subtype uint279_t is unsigned(278 downto 0);
constant uint279_t_SLV_LEN : integer := 279;
function uint279_t_to_slv(x : uint279_t) return std_logic_vector;
function slv_to_uint279_t(x : std_logic_vector) return uint279_t;
subtype int279_t is signed(278 downto 0);
constant int279_t_SLV_LEN : integer := 279;
function int279_t_to_slv(x : int279_t) return std_logic_vector;
function slv_to_int279_t(x : std_logic_vector) return int279_t;
subtype uint280_t is unsigned(279 downto 0);
constant uint280_t_SLV_LEN : integer := 280;
function uint280_t_to_slv(x : uint280_t) return std_logic_vector;
function slv_to_uint280_t(x : std_logic_vector) return uint280_t;
subtype int280_t is signed(279 downto 0);
constant int280_t_SLV_LEN : integer := 280;
function int280_t_to_slv(x : int280_t) return std_logic_vector;
function slv_to_int280_t(x : std_logic_vector) return int280_t;
subtype uint281_t is unsigned(280 downto 0);
constant uint281_t_SLV_LEN : integer := 281;
function uint281_t_to_slv(x : uint281_t) return std_logic_vector;
function slv_to_uint281_t(x : std_logic_vector) return uint281_t;
subtype int281_t is signed(280 downto 0);
constant int281_t_SLV_LEN : integer := 281;
function int281_t_to_slv(x : int281_t) return std_logic_vector;
function slv_to_int281_t(x : std_logic_vector) return int281_t;
subtype uint282_t is unsigned(281 downto 0);
constant uint282_t_SLV_LEN : integer := 282;
function uint282_t_to_slv(x : uint282_t) return std_logic_vector;
function slv_to_uint282_t(x : std_logic_vector) return uint282_t;
subtype int282_t is signed(281 downto 0);
constant int282_t_SLV_LEN : integer := 282;
function int282_t_to_slv(x : int282_t) return std_logic_vector;
function slv_to_int282_t(x : std_logic_vector) return int282_t;
subtype uint283_t is unsigned(282 downto 0);
constant uint283_t_SLV_LEN : integer := 283;
function uint283_t_to_slv(x : uint283_t) return std_logic_vector;
function slv_to_uint283_t(x : std_logic_vector) return uint283_t;
subtype int283_t is signed(282 downto 0);
constant int283_t_SLV_LEN : integer := 283;
function int283_t_to_slv(x : int283_t) return std_logic_vector;
function slv_to_int283_t(x : std_logic_vector) return int283_t;
subtype uint284_t is unsigned(283 downto 0);
constant uint284_t_SLV_LEN : integer := 284;
function uint284_t_to_slv(x : uint284_t) return std_logic_vector;
function slv_to_uint284_t(x : std_logic_vector) return uint284_t;
subtype int284_t is signed(283 downto 0);
constant int284_t_SLV_LEN : integer := 284;
function int284_t_to_slv(x : int284_t) return std_logic_vector;
function slv_to_int284_t(x : std_logic_vector) return int284_t;
subtype uint285_t is unsigned(284 downto 0);
constant uint285_t_SLV_LEN : integer := 285;
function uint285_t_to_slv(x : uint285_t) return std_logic_vector;
function slv_to_uint285_t(x : std_logic_vector) return uint285_t;
subtype int285_t is signed(284 downto 0);
constant int285_t_SLV_LEN : integer := 285;
function int285_t_to_slv(x : int285_t) return std_logic_vector;
function slv_to_int285_t(x : std_logic_vector) return int285_t;
subtype uint286_t is unsigned(285 downto 0);
constant uint286_t_SLV_LEN : integer := 286;
function uint286_t_to_slv(x : uint286_t) return std_logic_vector;
function slv_to_uint286_t(x : std_logic_vector) return uint286_t;
subtype int286_t is signed(285 downto 0);
constant int286_t_SLV_LEN : integer := 286;
function int286_t_to_slv(x : int286_t) return std_logic_vector;
function slv_to_int286_t(x : std_logic_vector) return int286_t;
subtype uint287_t is unsigned(286 downto 0);
constant uint287_t_SLV_LEN : integer := 287;
function uint287_t_to_slv(x : uint287_t) return std_logic_vector;
function slv_to_uint287_t(x : std_logic_vector) return uint287_t;
subtype int287_t is signed(286 downto 0);
constant int287_t_SLV_LEN : integer := 287;
function int287_t_to_slv(x : int287_t) return std_logic_vector;
function slv_to_int287_t(x : std_logic_vector) return int287_t;
subtype uint288_t is unsigned(287 downto 0);
constant uint288_t_SLV_LEN : integer := 288;
function uint288_t_to_slv(x : uint288_t) return std_logic_vector;
function slv_to_uint288_t(x : std_logic_vector) return uint288_t;
subtype int288_t is signed(287 downto 0);
constant int288_t_SLV_LEN : integer := 288;
function int288_t_to_slv(x : int288_t) return std_logic_vector;
function slv_to_int288_t(x : std_logic_vector) return int288_t;
subtype uint289_t is unsigned(288 downto 0);
constant uint289_t_SLV_LEN : integer := 289;
function uint289_t_to_slv(x : uint289_t) return std_logic_vector;
function slv_to_uint289_t(x : std_logic_vector) return uint289_t;
subtype int289_t is signed(288 downto 0);
constant int289_t_SLV_LEN : integer := 289;
function int289_t_to_slv(x : int289_t) return std_logic_vector;
function slv_to_int289_t(x : std_logic_vector) return int289_t;
subtype uint290_t is unsigned(289 downto 0);
constant uint290_t_SLV_LEN : integer := 290;
function uint290_t_to_slv(x : uint290_t) return std_logic_vector;
function slv_to_uint290_t(x : std_logic_vector) return uint290_t;
subtype int290_t is signed(289 downto 0);
constant int290_t_SLV_LEN : integer := 290;
function int290_t_to_slv(x : int290_t) return std_logic_vector;
function slv_to_int290_t(x : std_logic_vector) return int290_t;
subtype uint291_t is unsigned(290 downto 0);
constant uint291_t_SLV_LEN : integer := 291;
function uint291_t_to_slv(x : uint291_t) return std_logic_vector;
function slv_to_uint291_t(x : std_logic_vector) return uint291_t;
subtype int291_t is signed(290 downto 0);
constant int291_t_SLV_LEN : integer := 291;
function int291_t_to_slv(x : int291_t) return std_logic_vector;
function slv_to_int291_t(x : std_logic_vector) return int291_t;
subtype uint292_t is unsigned(291 downto 0);
constant uint292_t_SLV_LEN : integer := 292;
function uint292_t_to_slv(x : uint292_t) return std_logic_vector;
function slv_to_uint292_t(x : std_logic_vector) return uint292_t;
subtype int292_t is signed(291 downto 0);
constant int292_t_SLV_LEN : integer := 292;
function int292_t_to_slv(x : int292_t) return std_logic_vector;
function slv_to_int292_t(x : std_logic_vector) return int292_t;
subtype uint293_t is unsigned(292 downto 0);
constant uint293_t_SLV_LEN : integer := 293;
function uint293_t_to_slv(x : uint293_t) return std_logic_vector;
function slv_to_uint293_t(x : std_logic_vector) return uint293_t;
subtype int293_t is signed(292 downto 0);
constant int293_t_SLV_LEN : integer := 293;
function int293_t_to_slv(x : int293_t) return std_logic_vector;
function slv_to_int293_t(x : std_logic_vector) return int293_t;
subtype uint294_t is unsigned(293 downto 0);
constant uint294_t_SLV_LEN : integer := 294;
function uint294_t_to_slv(x : uint294_t) return std_logic_vector;
function slv_to_uint294_t(x : std_logic_vector) return uint294_t;
subtype int294_t is signed(293 downto 0);
constant int294_t_SLV_LEN : integer := 294;
function int294_t_to_slv(x : int294_t) return std_logic_vector;
function slv_to_int294_t(x : std_logic_vector) return int294_t;
subtype uint295_t is unsigned(294 downto 0);
constant uint295_t_SLV_LEN : integer := 295;
function uint295_t_to_slv(x : uint295_t) return std_logic_vector;
function slv_to_uint295_t(x : std_logic_vector) return uint295_t;
subtype int295_t is signed(294 downto 0);
constant int295_t_SLV_LEN : integer := 295;
function int295_t_to_slv(x : int295_t) return std_logic_vector;
function slv_to_int295_t(x : std_logic_vector) return int295_t;
subtype uint296_t is unsigned(295 downto 0);
constant uint296_t_SLV_LEN : integer := 296;
function uint296_t_to_slv(x : uint296_t) return std_logic_vector;
function slv_to_uint296_t(x : std_logic_vector) return uint296_t;
subtype int296_t is signed(295 downto 0);
constant int296_t_SLV_LEN : integer := 296;
function int296_t_to_slv(x : int296_t) return std_logic_vector;
function slv_to_int296_t(x : std_logic_vector) return int296_t;
subtype uint297_t is unsigned(296 downto 0);
constant uint297_t_SLV_LEN : integer := 297;
function uint297_t_to_slv(x : uint297_t) return std_logic_vector;
function slv_to_uint297_t(x : std_logic_vector) return uint297_t;
subtype int297_t is signed(296 downto 0);
constant int297_t_SLV_LEN : integer := 297;
function int297_t_to_slv(x : int297_t) return std_logic_vector;
function slv_to_int297_t(x : std_logic_vector) return int297_t;
subtype uint298_t is unsigned(297 downto 0);
constant uint298_t_SLV_LEN : integer := 298;
function uint298_t_to_slv(x : uint298_t) return std_logic_vector;
function slv_to_uint298_t(x : std_logic_vector) return uint298_t;
subtype int298_t is signed(297 downto 0);
constant int298_t_SLV_LEN : integer := 298;
function int298_t_to_slv(x : int298_t) return std_logic_vector;
function slv_to_int298_t(x : std_logic_vector) return int298_t;
subtype uint299_t is unsigned(298 downto 0);
constant uint299_t_SLV_LEN : integer := 299;
function uint299_t_to_slv(x : uint299_t) return std_logic_vector;
function slv_to_uint299_t(x : std_logic_vector) return uint299_t;
subtype int299_t is signed(298 downto 0);
constant int299_t_SLV_LEN : integer := 299;
function int299_t_to_slv(x : int299_t) return std_logic_vector;
function slv_to_int299_t(x : std_logic_vector) return int299_t;
subtype uint300_t is unsigned(299 downto 0);
constant uint300_t_SLV_LEN : integer := 300;
function uint300_t_to_slv(x : uint300_t) return std_logic_vector;
function slv_to_uint300_t(x : std_logic_vector) return uint300_t;
subtype int300_t is signed(299 downto 0);
constant int300_t_SLV_LEN : integer := 300;
function int300_t_to_slv(x : int300_t) return std_logic_vector;
function slv_to_int300_t(x : std_logic_vector) return int300_t;
subtype uint301_t is unsigned(300 downto 0);
constant uint301_t_SLV_LEN : integer := 301;
function uint301_t_to_slv(x : uint301_t) return std_logic_vector;
function slv_to_uint301_t(x : std_logic_vector) return uint301_t;
subtype int301_t is signed(300 downto 0);
constant int301_t_SLV_LEN : integer := 301;
function int301_t_to_slv(x : int301_t) return std_logic_vector;
function slv_to_int301_t(x : std_logic_vector) return int301_t;
subtype uint302_t is unsigned(301 downto 0);
constant uint302_t_SLV_LEN : integer := 302;
function uint302_t_to_slv(x : uint302_t) return std_logic_vector;
function slv_to_uint302_t(x : std_logic_vector) return uint302_t;
subtype int302_t is signed(301 downto 0);
constant int302_t_SLV_LEN : integer := 302;
function int302_t_to_slv(x : int302_t) return std_logic_vector;
function slv_to_int302_t(x : std_logic_vector) return int302_t;
subtype uint303_t is unsigned(302 downto 0);
constant uint303_t_SLV_LEN : integer := 303;
function uint303_t_to_slv(x : uint303_t) return std_logic_vector;
function slv_to_uint303_t(x : std_logic_vector) return uint303_t;
subtype int303_t is signed(302 downto 0);
constant int303_t_SLV_LEN : integer := 303;
function int303_t_to_slv(x : int303_t) return std_logic_vector;
function slv_to_int303_t(x : std_logic_vector) return int303_t;
subtype uint304_t is unsigned(303 downto 0);
constant uint304_t_SLV_LEN : integer := 304;
function uint304_t_to_slv(x : uint304_t) return std_logic_vector;
function slv_to_uint304_t(x : std_logic_vector) return uint304_t;
subtype int304_t is signed(303 downto 0);
constant int304_t_SLV_LEN : integer := 304;
function int304_t_to_slv(x : int304_t) return std_logic_vector;
function slv_to_int304_t(x : std_logic_vector) return int304_t;
subtype uint305_t is unsigned(304 downto 0);
constant uint305_t_SLV_LEN : integer := 305;
function uint305_t_to_slv(x : uint305_t) return std_logic_vector;
function slv_to_uint305_t(x : std_logic_vector) return uint305_t;
subtype int305_t is signed(304 downto 0);
constant int305_t_SLV_LEN : integer := 305;
function int305_t_to_slv(x : int305_t) return std_logic_vector;
function slv_to_int305_t(x : std_logic_vector) return int305_t;
subtype uint306_t is unsigned(305 downto 0);
constant uint306_t_SLV_LEN : integer := 306;
function uint306_t_to_slv(x : uint306_t) return std_logic_vector;
function slv_to_uint306_t(x : std_logic_vector) return uint306_t;
subtype int306_t is signed(305 downto 0);
constant int306_t_SLV_LEN : integer := 306;
function int306_t_to_slv(x : int306_t) return std_logic_vector;
function slv_to_int306_t(x : std_logic_vector) return int306_t;
subtype uint307_t is unsigned(306 downto 0);
constant uint307_t_SLV_LEN : integer := 307;
function uint307_t_to_slv(x : uint307_t) return std_logic_vector;
function slv_to_uint307_t(x : std_logic_vector) return uint307_t;
subtype int307_t is signed(306 downto 0);
constant int307_t_SLV_LEN : integer := 307;
function int307_t_to_slv(x : int307_t) return std_logic_vector;
function slv_to_int307_t(x : std_logic_vector) return int307_t;
subtype uint308_t is unsigned(307 downto 0);
constant uint308_t_SLV_LEN : integer := 308;
function uint308_t_to_slv(x : uint308_t) return std_logic_vector;
function slv_to_uint308_t(x : std_logic_vector) return uint308_t;
subtype int308_t is signed(307 downto 0);
constant int308_t_SLV_LEN : integer := 308;
function int308_t_to_slv(x : int308_t) return std_logic_vector;
function slv_to_int308_t(x : std_logic_vector) return int308_t;
subtype uint309_t is unsigned(308 downto 0);
constant uint309_t_SLV_LEN : integer := 309;
function uint309_t_to_slv(x : uint309_t) return std_logic_vector;
function slv_to_uint309_t(x : std_logic_vector) return uint309_t;
subtype int309_t is signed(308 downto 0);
constant int309_t_SLV_LEN : integer := 309;
function int309_t_to_slv(x : int309_t) return std_logic_vector;
function slv_to_int309_t(x : std_logic_vector) return int309_t;
subtype uint310_t is unsigned(309 downto 0);
constant uint310_t_SLV_LEN : integer := 310;
function uint310_t_to_slv(x : uint310_t) return std_logic_vector;
function slv_to_uint310_t(x : std_logic_vector) return uint310_t;
subtype int310_t is signed(309 downto 0);
constant int310_t_SLV_LEN : integer := 310;
function int310_t_to_slv(x : int310_t) return std_logic_vector;
function slv_to_int310_t(x : std_logic_vector) return int310_t;
subtype uint311_t is unsigned(310 downto 0);
constant uint311_t_SLV_LEN : integer := 311;
function uint311_t_to_slv(x : uint311_t) return std_logic_vector;
function slv_to_uint311_t(x : std_logic_vector) return uint311_t;
subtype int311_t is signed(310 downto 0);
constant int311_t_SLV_LEN : integer := 311;
function int311_t_to_slv(x : int311_t) return std_logic_vector;
function slv_to_int311_t(x : std_logic_vector) return int311_t;
subtype uint312_t is unsigned(311 downto 0);
constant uint312_t_SLV_LEN : integer := 312;
function uint312_t_to_slv(x : uint312_t) return std_logic_vector;
function slv_to_uint312_t(x : std_logic_vector) return uint312_t;
subtype int312_t is signed(311 downto 0);
constant int312_t_SLV_LEN : integer := 312;
function int312_t_to_slv(x : int312_t) return std_logic_vector;
function slv_to_int312_t(x : std_logic_vector) return int312_t;
subtype uint313_t is unsigned(312 downto 0);
constant uint313_t_SLV_LEN : integer := 313;
function uint313_t_to_slv(x : uint313_t) return std_logic_vector;
function slv_to_uint313_t(x : std_logic_vector) return uint313_t;
subtype int313_t is signed(312 downto 0);
constant int313_t_SLV_LEN : integer := 313;
function int313_t_to_slv(x : int313_t) return std_logic_vector;
function slv_to_int313_t(x : std_logic_vector) return int313_t;
subtype uint314_t is unsigned(313 downto 0);
constant uint314_t_SLV_LEN : integer := 314;
function uint314_t_to_slv(x : uint314_t) return std_logic_vector;
function slv_to_uint314_t(x : std_logic_vector) return uint314_t;
subtype int314_t is signed(313 downto 0);
constant int314_t_SLV_LEN : integer := 314;
function int314_t_to_slv(x : int314_t) return std_logic_vector;
function slv_to_int314_t(x : std_logic_vector) return int314_t;
subtype uint315_t is unsigned(314 downto 0);
constant uint315_t_SLV_LEN : integer := 315;
function uint315_t_to_slv(x : uint315_t) return std_logic_vector;
function slv_to_uint315_t(x : std_logic_vector) return uint315_t;
subtype int315_t is signed(314 downto 0);
constant int315_t_SLV_LEN : integer := 315;
function int315_t_to_slv(x : int315_t) return std_logic_vector;
function slv_to_int315_t(x : std_logic_vector) return int315_t;
subtype uint316_t is unsigned(315 downto 0);
constant uint316_t_SLV_LEN : integer := 316;
function uint316_t_to_slv(x : uint316_t) return std_logic_vector;
function slv_to_uint316_t(x : std_logic_vector) return uint316_t;
subtype int316_t is signed(315 downto 0);
constant int316_t_SLV_LEN : integer := 316;
function int316_t_to_slv(x : int316_t) return std_logic_vector;
function slv_to_int316_t(x : std_logic_vector) return int316_t;
subtype uint317_t is unsigned(316 downto 0);
constant uint317_t_SLV_LEN : integer := 317;
function uint317_t_to_slv(x : uint317_t) return std_logic_vector;
function slv_to_uint317_t(x : std_logic_vector) return uint317_t;
subtype int317_t is signed(316 downto 0);
constant int317_t_SLV_LEN : integer := 317;
function int317_t_to_slv(x : int317_t) return std_logic_vector;
function slv_to_int317_t(x : std_logic_vector) return int317_t;
subtype uint318_t is unsigned(317 downto 0);
constant uint318_t_SLV_LEN : integer := 318;
function uint318_t_to_slv(x : uint318_t) return std_logic_vector;
function slv_to_uint318_t(x : std_logic_vector) return uint318_t;
subtype int318_t is signed(317 downto 0);
constant int318_t_SLV_LEN : integer := 318;
function int318_t_to_slv(x : int318_t) return std_logic_vector;
function slv_to_int318_t(x : std_logic_vector) return int318_t;
subtype uint319_t is unsigned(318 downto 0);
constant uint319_t_SLV_LEN : integer := 319;
function uint319_t_to_slv(x : uint319_t) return std_logic_vector;
function slv_to_uint319_t(x : std_logic_vector) return uint319_t;
subtype int319_t is signed(318 downto 0);
constant int319_t_SLV_LEN : integer := 319;
function int319_t_to_slv(x : int319_t) return std_logic_vector;
function slv_to_int319_t(x : std_logic_vector) return int319_t;
subtype uint320_t is unsigned(319 downto 0);
constant uint320_t_SLV_LEN : integer := 320;
function uint320_t_to_slv(x : uint320_t) return std_logic_vector;
function slv_to_uint320_t(x : std_logic_vector) return uint320_t;
subtype int320_t is signed(319 downto 0);
constant int320_t_SLV_LEN : integer := 320;
function int320_t_to_slv(x : int320_t) return std_logic_vector;
function slv_to_int320_t(x : std_logic_vector) return int320_t;
subtype uint321_t is unsigned(320 downto 0);
constant uint321_t_SLV_LEN : integer := 321;
function uint321_t_to_slv(x : uint321_t) return std_logic_vector;
function slv_to_uint321_t(x : std_logic_vector) return uint321_t;
subtype int321_t is signed(320 downto 0);
constant int321_t_SLV_LEN : integer := 321;
function int321_t_to_slv(x : int321_t) return std_logic_vector;
function slv_to_int321_t(x : std_logic_vector) return int321_t;
subtype uint322_t is unsigned(321 downto 0);
constant uint322_t_SLV_LEN : integer := 322;
function uint322_t_to_slv(x : uint322_t) return std_logic_vector;
function slv_to_uint322_t(x : std_logic_vector) return uint322_t;
subtype int322_t is signed(321 downto 0);
constant int322_t_SLV_LEN : integer := 322;
function int322_t_to_slv(x : int322_t) return std_logic_vector;
function slv_to_int322_t(x : std_logic_vector) return int322_t;
subtype uint323_t is unsigned(322 downto 0);
constant uint323_t_SLV_LEN : integer := 323;
function uint323_t_to_slv(x : uint323_t) return std_logic_vector;
function slv_to_uint323_t(x : std_logic_vector) return uint323_t;
subtype int323_t is signed(322 downto 0);
constant int323_t_SLV_LEN : integer := 323;
function int323_t_to_slv(x : int323_t) return std_logic_vector;
function slv_to_int323_t(x : std_logic_vector) return int323_t;
subtype uint324_t is unsigned(323 downto 0);
constant uint324_t_SLV_LEN : integer := 324;
function uint324_t_to_slv(x : uint324_t) return std_logic_vector;
function slv_to_uint324_t(x : std_logic_vector) return uint324_t;
subtype int324_t is signed(323 downto 0);
constant int324_t_SLV_LEN : integer := 324;
function int324_t_to_slv(x : int324_t) return std_logic_vector;
function slv_to_int324_t(x : std_logic_vector) return int324_t;
subtype uint325_t is unsigned(324 downto 0);
constant uint325_t_SLV_LEN : integer := 325;
function uint325_t_to_slv(x : uint325_t) return std_logic_vector;
function slv_to_uint325_t(x : std_logic_vector) return uint325_t;
subtype int325_t is signed(324 downto 0);
constant int325_t_SLV_LEN : integer := 325;
function int325_t_to_slv(x : int325_t) return std_logic_vector;
function slv_to_int325_t(x : std_logic_vector) return int325_t;
subtype uint326_t is unsigned(325 downto 0);
constant uint326_t_SLV_LEN : integer := 326;
function uint326_t_to_slv(x : uint326_t) return std_logic_vector;
function slv_to_uint326_t(x : std_logic_vector) return uint326_t;
subtype int326_t is signed(325 downto 0);
constant int326_t_SLV_LEN : integer := 326;
function int326_t_to_slv(x : int326_t) return std_logic_vector;
function slv_to_int326_t(x : std_logic_vector) return int326_t;
subtype uint327_t is unsigned(326 downto 0);
constant uint327_t_SLV_LEN : integer := 327;
function uint327_t_to_slv(x : uint327_t) return std_logic_vector;
function slv_to_uint327_t(x : std_logic_vector) return uint327_t;
subtype int327_t is signed(326 downto 0);
constant int327_t_SLV_LEN : integer := 327;
function int327_t_to_slv(x : int327_t) return std_logic_vector;
function slv_to_int327_t(x : std_logic_vector) return int327_t;
subtype uint328_t is unsigned(327 downto 0);
constant uint328_t_SLV_LEN : integer := 328;
function uint328_t_to_slv(x : uint328_t) return std_logic_vector;
function slv_to_uint328_t(x : std_logic_vector) return uint328_t;
subtype int328_t is signed(327 downto 0);
constant int328_t_SLV_LEN : integer := 328;
function int328_t_to_slv(x : int328_t) return std_logic_vector;
function slv_to_int328_t(x : std_logic_vector) return int328_t;
subtype uint329_t is unsigned(328 downto 0);
constant uint329_t_SLV_LEN : integer := 329;
function uint329_t_to_slv(x : uint329_t) return std_logic_vector;
function slv_to_uint329_t(x : std_logic_vector) return uint329_t;
subtype int329_t is signed(328 downto 0);
constant int329_t_SLV_LEN : integer := 329;
function int329_t_to_slv(x : int329_t) return std_logic_vector;
function slv_to_int329_t(x : std_logic_vector) return int329_t;
subtype uint330_t is unsigned(329 downto 0);
constant uint330_t_SLV_LEN : integer := 330;
function uint330_t_to_slv(x : uint330_t) return std_logic_vector;
function slv_to_uint330_t(x : std_logic_vector) return uint330_t;
subtype int330_t is signed(329 downto 0);
constant int330_t_SLV_LEN : integer := 330;
function int330_t_to_slv(x : int330_t) return std_logic_vector;
function slv_to_int330_t(x : std_logic_vector) return int330_t;
subtype uint331_t is unsigned(330 downto 0);
constant uint331_t_SLV_LEN : integer := 331;
function uint331_t_to_slv(x : uint331_t) return std_logic_vector;
function slv_to_uint331_t(x : std_logic_vector) return uint331_t;
subtype int331_t is signed(330 downto 0);
constant int331_t_SLV_LEN : integer := 331;
function int331_t_to_slv(x : int331_t) return std_logic_vector;
function slv_to_int331_t(x : std_logic_vector) return int331_t;
subtype uint332_t is unsigned(331 downto 0);
constant uint332_t_SLV_LEN : integer := 332;
function uint332_t_to_slv(x : uint332_t) return std_logic_vector;
function slv_to_uint332_t(x : std_logic_vector) return uint332_t;
subtype int332_t is signed(331 downto 0);
constant int332_t_SLV_LEN : integer := 332;
function int332_t_to_slv(x : int332_t) return std_logic_vector;
function slv_to_int332_t(x : std_logic_vector) return int332_t;
subtype uint333_t is unsigned(332 downto 0);
constant uint333_t_SLV_LEN : integer := 333;
function uint333_t_to_slv(x : uint333_t) return std_logic_vector;
function slv_to_uint333_t(x : std_logic_vector) return uint333_t;
subtype int333_t is signed(332 downto 0);
constant int333_t_SLV_LEN : integer := 333;
function int333_t_to_slv(x : int333_t) return std_logic_vector;
function slv_to_int333_t(x : std_logic_vector) return int333_t;
subtype uint334_t is unsigned(333 downto 0);
constant uint334_t_SLV_LEN : integer := 334;
function uint334_t_to_slv(x : uint334_t) return std_logic_vector;
function slv_to_uint334_t(x : std_logic_vector) return uint334_t;
subtype int334_t is signed(333 downto 0);
constant int334_t_SLV_LEN : integer := 334;
function int334_t_to_slv(x : int334_t) return std_logic_vector;
function slv_to_int334_t(x : std_logic_vector) return int334_t;
subtype uint335_t is unsigned(334 downto 0);
constant uint335_t_SLV_LEN : integer := 335;
function uint335_t_to_slv(x : uint335_t) return std_logic_vector;
function slv_to_uint335_t(x : std_logic_vector) return uint335_t;
subtype int335_t is signed(334 downto 0);
constant int335_t_SLV_LEN : integer := 335;
function int335_t_to_slv(x : int335_t) return std_logic_vector;
function slv_to_int335_t(x : std_logic_vector) return int335_t;
subtype uint336_t is unsigned(335 downto 0);
constant uint336_t_SLV_LEN : integer := 336;
function uint336_t_to_slv(x : uint336_t) return std_logic_vector;
function slv_to_uint336_t(x : std_logic_vector) return uint336_t;
subtype int336_t is signed(335 downto 0);
constant int336_t_SLV_LEN : integer := 336;
function int336_t_to_slv(x : int336_t) return std_logic_vector;
function slv_to_int336_t(x : std_logic_vector) return int336_t;
subtype uint337_t is unsigned(336 downto 0);
constant uint337_t_SLV_LEN : integer := 337;
function uint337_t_to_slv(x : uint337_t) return std_logic_vector;
function slv_to_uint337_t(x : std_logic_vector) return uint337_t;
subtype int337_t is signed(336 downto 0);
constant int337_t_SLV_LEN : integer := 337;
function int337_t_to_slv(x : int337_t) return std_logic_vector;
function slv_to_int337_t(x : std_logic_vector) return int337_t;
subtype uint338_t is unsigned(337 downto 0);
constant uint338_t_SLV_LEN : integer := 338;
function uint338_t_to_slv(x : uint338_t) return std_logic_vector;
function slv_to_uint338_t(x : std_logic_vector) return uint338_t;
subtype int338_t is signed(337 downto 0);
constant int338_t_SLV_LEN : integer := 338;
function int338_t_to_slv(x : int338_t) return std_logic_vector;
function slv_to_int338_t(x : std_logic_vector) return int338_t;
subtype uint339_t is unsigned(338 downto 0);
constant uint339_t_SLV_LEN : integer := 339;
function uint339_t_to_slv(x : uint339_t) return std_logic_vector;
function slv_to_uint339_t(x : std_logic_vector) return uint339_t;
subtype int339_t is signed(338 downto 0);
constant int339_t_SLV_LEN : integer := 339;
function int339_t_to_slv(x : int339_t) return std_logic_vector;
function slv_to_int339_t(x : std_logic_vector) return int339_t;
subtype uint340_t is unsigned(339 downto 0);
constant uint340_t_SLV_LEN : integer := 340;
function uint340_t_to_slv(x : uint340_t) return std_logic_vector;
function slv_to_uint340_t(x : std_logic_vector) return uint340_t;
subtype int340_t is signed(339 downto 0);
constant int340_t_SLV_LEN : integer := 340;
function int340_t_to_slv(x : int340_t) return std_logic_vector;
function slv_to_int340_t(x : std_logic_vector) return int340_t;
subtype uint341_t is unsigned(340 downto 0);
constant uint341_t_SLV_LEN : integer := 341;
function uint341_t_to_slv(x : uint341_t) return std_logic_vector;
function slv_to_uint341_t(x : std_logic_vector) return uint341_t;
subtype int341_t is signed(340 downto 0);
constant int341_t_SLV_LEN : integer := 341;
function int341_t_to_slv(x : int341_t) return std_logic_vector;
function slv_to_int341_t(x : std_logic_vector) return int341_t;
subtype uint342_t is unsigned(341 downto 0);
constant uint342_t_SLV_LEN : integer := 342;
function uint342_t_to_slv(x : uint342_t) return std_logic_vector;
function slv_to_uint342_t(x : std_logic_vector) return uint342_t;
subtype int342_t is signed(341 downto 0);
constant int342_t_SLV_LEN : integer := 342;
function int342_t_to_slv(x : int342_t) return std_logic_vector;
function slv_to_int342_t(x : std_logic_vector) return int342_t;
subtype uint343_t is unsigned(342 downto 0);
constant uint343_t_SLV_LEN : integer := 343;
function uint343_t_to_slv(x : uint343_t) return std_logic_vector;
function slv_to_uint343_t(x : std_logic_vector) return uint343_t;
subtype int343_t is signed(342 downto 0);
constant int343_t_SLV_LEN : integer := 343;
function int343_t_to_slv(x : int343_t) return std_logic_vector;
function slv_to_int343_t(x : std_logic_vector) return int343_t;
subtype uint344_t is unsigned(343 downto 0);
constant uint344_t_SLV_LEN : integer := 344;
function uint344_t_to_slv(x : uint344_t) return std_logic_vector;
function slv_to_uint344_t(x : std_logic_vector) return uint344_t;
subtype int344_t is signed(343 downto 0);
constant int344_t_SLV_LEN : integer := 344;
function int344_t_to_slv(x : int344_t) return std_logic_vector;
function slv_to_int344_t(x : std_logic_vector) return int344_t;
subtype uint345_t is unsigned(344 downto 0);
constant uint345_t_SLV_LEN : integer := 345;
function uint345_t_to_slv(x : uint345_t) return std_logic_vector;
function slv_to_uint345_t(x : std_logic_vector) return uint345_t;
subtype int345_t is signed(344 downto 0);
constant int345_t_SLV_LEN : integer := 345;
function int345_t_to_slv(x : int345_t) return std_logic_vector;
function slv_to_int345_t(x : std_logic_vector) return int345_t;
subtype uint346_t is unsigned(345 downto 0);
constant uint346_t_SLV_LEN : integer := 346;
function uint346_t_to_slv(x : uint346_t) return std_logic_vector;
function slv_to_uint346_t(x : std_logic_vector) return uint346_t;
subtype int346_t is signed(345 downto 0);
constant int346_t_SLV_LEN : integer := 346;
function int346_t_to_slv(x : int346_t) return std_logic_vector;
function slv_to_int346_t(x : std_logic_vector) return int346_t;
subtype uint347_t is unsigned(346 downto 0);
constant uint347_t_SLV_LEN : integer := 347;
function uint347_t_to_slv(x : uint347_t) return std_logic_vector;
function slv_to_uint347_t(x : std_logic_vector) return uint347_t;
subtype int347_t is signed(346 downto 0);
constant int347_t_SLV_LEN : integer := 347;
function int347_t_to_slv(x : int347_t) return std_logic_vector;
function slv_to_int347_t(x : std_logic_vector) return int347_t;
subtype uint348_t is unsigned(347 downto 0);
constant uint348_t_SLV_LEN : integer := 348;
function uint348_t_to_slv(x : uint348_t) return std_logic_vector;
function slv_to_uint348_t(x : std_logic_vector) return uint348_t;
subtype int348_t is signed(347 downto 0);
constant int348_t_SLV_LEN : integer := 348;
function int348_t_to_slv(x : int348_t) return std_logic_vector;
function slv_to_int348_t(x : std_logic_vector) return int348_t;
subtype uint349_t is unsigned(348 downto 0);
constant uint349_t_SLV_LEN : integer := 349;
function uint349_t_to_slv(x : uint349_t) return std_logic_vector;
function slv_to_uint349_t(x : std_logic_vector) return uint349_t;
subtype int349_t is signed(348 downto 0);
constant int349_t_SLV_LEN : integer := 349;
function int349_t_to_slv(x : int349_t) return std_logic_vector;
function slv_to_int349_t(x : std_logic_vector) return int349_t;
subtype uint350_t is unsigned(349 downto 0);
constant uint350_t_SLV_LEN : integer := 350;
function uint350_t_to_slv(x : uint350_t) return std_logic_vector;
function slv_to_uint350_t(x : std_logic_vector) return uint350_t;
subtype int350_t is signed(349 downto 0);
constant int350_t_SLV_LEN : integer := 350;
function int350_t_to_slv(x : int350_t) return std_logic_vector;
function slv_to_int350_t(x : std_logic_vector) return int350_t;
subtype uint351_t is unsigned(350 downto 0);
constant uint351_t_SLV_LEN : integer := 351;
function uint351_t_to_slv(x : uint351_t) return std_logic_vector;
function slv_to_uint351_t(x : std_logic_vector) return uint351_t;
subtype int351_t is signed(350 downto 0);
constant int351_t_SLV_LEN : integer := 351;
function int351_t_to_slv(x : int351_t) return std_logic_vector;
function slv_to_int351_t(x : std_logic_vector) return int351_t;
subtype uint352_t is unsigned(351 downto 0);
constant uint352_t_SLV_LEN : integer := 352;
function uint352_t_to_slv(x : uint352_t) return std_logic_vector;
function slv_to_uint352_t(x : std_logic_vector) return uint352_t;
subtype int352_t is signed(351 downto 0);
constant int352_t_SLV_LEN : integer := 352;
function int352_t_to_slv(x : int352_t) return std_logic_vector;
function slv_to_int352_t(x : std_logic_vector) return int352_t;
subtype uint353_t is unsigned(352 downto 0);
constant uint353_t_SLV_LEN : integer := 353;
function uint353_t_to_slv(x : uint353_t) return std_logic_vector;
function slv_to_uint353_t(x : std_logic_vector) return uint353_t;
subtype int353_t is signed(352 downto 0);
constant int353_t_SLV_LEN : integer := 353;
function int353_t_to_slv(x : int353_t) return std_logic_vector;
function slv_to_int353_t(x : std_logic_vector) return int353_t;
subtype uint354_t is unsigned(353 downto 0);
constant uint354_t_SLV_LEN : integer := 354;
function uint354_t_to_slv(x : uint354_t) return std_logic_vector;
function slv_to_uint354_t(x : std_logic_vector) return uint354_t;
subtype int354_t is signed(353 downto 0);
constant int354_t_SLV_LEN : integer := 354;
function int354_t_to_slv(x : int354_t) return std_logic_vector;
function slv_to_int354_t(x : std_logic_vector) return int354_t;
subtype uint355_t is unsigned(354 downto 0);
constant uint355_t_SLV_LEN : integer := 355;
function uint355_t_to_slv(x : uint355_t) return std_logic_vector;
function slv_to_uint355_t(x : std_logic_vector) return uint355_t;
subtype int355_t is signed(354 downto 0);
constant int355_t_SLV_LEN : integer := 355;
function int355_t_to_slv(x : int355_t) return std_logic_vector;
function slv_to_int355_t(x : std_logic_vector) return int355_t;
subtype uint356_t is unsigned(355 downto 0);
constant uint356_t_SLV_LEN : integer := 356;
function uint356_t_to_slv(x : uint356_t) return std_logic_vector;
function slv_to_uint356_t(x : std_logic_vector) return uint356_t;
subtype int356_t is signed(355 downto 0);
constant int356_t_SLV_LEN : integer := 356;
function int356_t_to_slv(x : int356_t) return std_logic_vector;
function slv_to_int356_t(x : std_logic_vector) return int356_t;
subtype uint357_t is unsigned(356 downto 0);
constant uint357_t_SLV_LEN : integer := 357;
function uint357_t_to_slv(x : uint357_t) return std_logic_vector;
function slv_to_uint357_t(x : std_logic_vector) return uint357_t;
subtype int357_t is signed(356 downto 0);
constant int357_t_SLV_LEN : integer := 357;
function int357_t_to_slv(x : int357_t) return std_logic_vector;
function slv_to_int357_t(x : std_logic_vector) return int357_t;
subtype uint358_t is unsigned(357 downto 0);
constant uint358_t_SLV_LEN : integer := 358;
function uint358_t_to_slv(x : uint358_t) return std_logic_vector;
function slv_to_uint358_t(x : std_logic_vector) return uint358_t;
subtype int358_t is signed(357 downto 0);
constant int358_t_SLV_LEN : integer := 358;
function int358_t_to_slv(x : int358_t) return std_logic_vector;
function slv_to_int358_t(x : std_logic_vector) return int358_t;
subtype uint359_t is unsigned(358 downto 0);
constant uint359_t_SLV_LEN : integer := 359;
function uint359_t_to_slv(x : uint359_t) return std_logic_vector;
function slv_to_uint359_t(x : std_logic_vector) return uint359_t;
subtype int359_t is signed(358 downto 0);
constant int359_t_SLV_LEN : integer := 359;
function int359_t_to_slv(x : int359_t) return std_logic_vector;
function slv_to_int359_t(x : std_logic_vector) return int359_t;
subtype uint360_t is unsigned(359 downto 0);
constant uint360_t_SLV_LEN : integer := 360;
function uint360_t_to_slv(x : uint360_t) return std_logic_vector;
function slv_to_uint360_t(x : std_logic_vector) return uint360_t;
subtype int360_t is signed(359 downto 0);
constant int360_t_SLV_LEN : integer := 360;
function int360_t_to_slv(x : int360_t) return std_logic_vector;
function slv_to_int360_t(x : std_logic_vector) return int360_t;
subtype uint361_t is unsigned(360 downto 0);
constant uint361_t_SLV_LEN : integer := 361;
function uint361_t_to_slv(x : uint361_t) return std_logic_vector;
function slv_to_uint361_t(x : std_logic_vector) return uint361_t;
subtype int361_t is signed(360 downto 0);
constant int361_t_SLV_LEN : integer := 361;
function int361_t_to_slv(x : int361_t) return std_logic_vector;
function slv_to_int361_t(x : std_logic_vector) return int361_t;
subtype uint362_t is unsigned(361 downto 0);
constant uint362_t_SLV_LEN : integer := 362;
function uint362_t_to_slv(x : uint362_t) return std_logic_vector;
function slv_to_uint362_t(x : std_logic_vector) return uint362_t;
subtype int362_t is signed(361 downto 0);
constant int362_t_SLV_LEN : integer := 362;
function int362_t_to_slv(x : int362_t) return std_logic_vector;
function slv_to_int362_t(x : std_logic_vector) return int362_t;
subtype uint363_t is unsigned(362 downto 0);
constant uint363_t_SLV_LEN : integer := 363;
function uint363_t_to_slv(x : uint363_t) return std_logic_vector;
function slv_to_uint363_t(x : std_logic_vector) return uint363_t;
subtype int363_t is signed(362 downto 0);
constant int363_t_SLV_LEN : integer := 363;
function int363_t_to_slv(x : int363_t) return std_logic_vector;
function slv_to_int363_t(x : std_logic_vector) return int363_t;
subtype uint364_t is unsigned(363 downto 0);
constant uint364_t_SLV_LEN : integer := 364;
function uint364_t_to_slv(x : uint364_t) return std_logic_vector;
function slv_to_uint364_t(x : std_logic_vector) return uint364_t;
subtype int364_t is signed(363 downto 0);
constant int364_t_SLV_LEN : integer := 364;
function int364_t_to_slv(x : int364_t) return std_logic_vector;
function slv_to_int364_t(x : std_logic_vector) return int364_t;
subtype uint365_t is unsigned(364 downto 0);
constant uint365_t_SLV_LEN : integer := 365;
function uint365_t_to_slv(x : uint365_t) return std_logic_vector;
function slv_to_uint365_t(x : std_logic_vector) return uint365_t;
subtype int365_t is signed(364 downto 0);
constant int365_t_SLV_LEN : integer := 365;
function int365_t_to_slv(x : int365_t) return std_logic_vector;
function slv_to_int365_t(x : std_logic_vector) return int365_t;
subtype uint366_t is unsigned(365 downto 0);
constant uint366_t_SLV_LEN : integer := 366;
function uint366_t_to_slv(x : uint366_t) return std_logic_vector;
function slv_to_uint366_t(x : std_logic_vector) return uint366_t;
subtype int366_t is signed(365 downto 0);
constant int366_t_SLV_LEN : integer := 366;
function int366_t_to_slv(x : int366_t) return std_logic_vector;
function slv_to_int366_t(x : std_logic_vector) return int366_t;
subtype uint367_t is unsigned(366 downto 0);
constant uint367_t_SLV_LEN : integer := 367;
function uint367_t_to_slv(x : uint367_t) return std_logic_vector;
function slv_to_uint367_t(x : std_logic_vector) return uint367_t;
subtype int367_t is signed(366 downto 0);
constant int367_t_SLV_LEN : integer := 367;
function int367_t_to_slv(x : int367_t) return std_logic_vector;
function slv_to_int367_t(x : std_logic_vector) return int367_t;
subtype uint368_t is unsigned(367 downto 0);
constant uint368_t_SLV_LEN : integer := 368;
function uint368_t_to_slv(x : uint368_t) return std_logic_vector;
function slv_to_uint368_t(x : std_logic_vector) return uint368_t;
subtype int368_t is signed(367 downto 0);
constant int368_t_SLV_LEN : integer := 368;
function int368_t_to_slv(x : int368_t) return std_logic_vector;
function slv_to_int368_t(x : std_logic_vector) return int368_t;
subtype uint369_t is unsigned(368 downto 0);
constant uint369_t_SLV_LEN : integer := 369;
function uint369_t_to_slv(x : uint369_t) return std_logic_vector;
function slv_to_uint369_t(x : std_logic_vector) return uint369_t;
subtype int369_t is signed(368 downto 0);
constant int369_t_SLV_LEN : integer := 369;
function int369_t_to_slv(x : int369_t) return std_logic_vector;
function slv_to_int369_t(x : std_logic_vector) return int369_t;
subtype uint370_t is unsigned(369 downto 0);
constant uint370_t_SLV_LEN : integer := 370;
function uint370_t_to_slv(x : uint370_t) return std_logic_vector;
function slv_to_uint370_t(x : std_logic_vector) return uint370_t;
subtype int370_t is signed(369 downto 0);
constant int370_t_SLV_LEN : integer := 370;
function int370_t_to_slv(x : int370_t) return std_logic_vector;
function slv_to_int370_t(x : std_logic_vector) return int370_t;
subtype uint371_t is unsigned(370 downto 0);
constant uint371_t_SLV_LEN : integer := 371;
function uint371_t_to_slv(x : uint371_t) return std_logic_vector;
function slv_to_uint371_t(x : std_logic_vector) return uint371_t;
subtype int371_t is signed(370 downto 0);
constant int371_t_SLV_LEN : integer := 371;
function int371_t_to_slv(x : int371_t) return std_logic_vector;
function slv_to_int371_t(x : std_logic_vector) return int371_t;
subtype uint372_t is unsigned(371 downto 0);
constant uint372_t_SLV_LEN : integer := 372;
function uint372_t_to_slv(x : uint372_t) return std_logic_vector;
function slv_to_uint372_t(x : std_logic_vector) return uint372_t;
subtype int372_t is signed(371 downto 0);
constant int372_t_SLV_LEN : integer := 372;
function int372_t_to_slv(x : int372_t) return std_logic_vector;
function slv_to_int372_t(x : std_logic_vector) return int372_t;
subtype uint373_t is unsigned(372 downto 0);
constant uint373_t_SLV_LEN : integer := 373;
function uint373_t_to_slv(x : uint373_t) return std_logic_vector;
function slv_to_uint373_t(x : std_logic_vector) return uint373_t;
subtype int373_t is signed(372 downto 0);
constant int373_t_SLV_LEN : integer := 373;
function int373_t_to_slv(x : int373_t) return std_logic_vector;
function slv_to_int373_t(x : std_logic_vector) return int373_t;
subtype uint374_t is unsigned(373 downto 0);
constant uint374_t_SLV_LEN : integer := 374;
function uint374_t_to_slv(x : uint374_t) return std_logic_vector;
function slv_to_uint374_t(x : std_logic_vector) return uint374_t;
subtype int374_t is signed(373 downto 0);
constant int374_t_SLV_LEN : integer := 374;
function int374_t_to_slv(x : int374_t) return std_logic_vector;
function slv_to_int374_t(x : std_logic_vector) return int374_t;
subtype uint375_t is unsigned(374 downto 0);
constant uint375_t_SLV_LEN : integer := 375;
function uint375_t_to_slv(x : uint375_t) return std_logic_vector;
function slv_to_uint375_t(x : std_logic_vector) return uint375_t;
subtype int375_t is signed(374 downto 0);
constant int375_t_SLV_LEN : integer := 375;
function int375_t_to_slv(x : int375_t) return std_logic_vector;
function slv_to_int375_t(x : std_logic_vector) return int375_t;
subtype uint376_t is unsigned(375 downto 0);
constant uint376_t_SLV_LEN : integer := 376;
function uint376_t_to_slv(x : uint376_t) return std_logic_vector;
function slv_to_uint376_t(x : std_logic_vector) return uint376_t;
subtype int376_t is signed(375 downto 0);
constant int376_t_SLV_LEN : integer := 376;
function int376_t_to_slv(x : int376_t) return std_logic_vector;
function slv_to_int376_t(x : std_logic_vector) return int376_t;
subtype uint377_t is unsigned(376 downto 0);
constant uint377_t_SLV_LEN : integer := 377;
function uint377_t_to_slv(x : uint377_t) return std_logic_vector;
function slv_to_uint377_t(x : std_logic_vector) return uint377_t;
subtype int377_t is signed(376 downto 0);
constant int377_t_SLV_LEN : integer := 377;
function int377_t_to_slv(x : int377_t) return std_logic_vector;
function slv_to_int377_t(x : std_logic_vector) return int377_t;
subtype uint378_t is unsigned(377 downto 0);
constant uint378_t_SLV_LEN : integer := 378;
function uint378_t_to_slv(x : uint378_t) return std_logic_vector;
function slv_to_uint378_t(x : std_logic_vector) return uint378_t;
subtype int378_t is signed(377 downto 0);
constant int378_t_SLV_LEN : integer := 378;
function int378_t_to_slv(x : int378_t) return std_logic_vector;
function slv_to_int378_t(x : std_logic_vector) return int378_t;
subtype uint379_t is unsigned(378 downto 0);
constant uint379_t_SLV_LEN : integer := 379;
function uint379_t_to_slv(x : uint379_t) return std_logic_vector;
function slv_to_uint379_t(x : std_logic_vector) return uint379_t;
subtype int379_t is signed(378 downto 0);
constant int379_t_SLV_LEN : integer := 379;
function int379_t_to_slv(x : int379_t) return std_logic_vector;
function slv_to_int379_t(x : std_logic_vector) return int379_t;
subtype uint380_t is unsigned(379 downto 0);
constant uint380_t_SLV_LEN : integer := 380;
function uint380_t_to_slv(x : uint380_t) return std_logic_vector;
function slv_to_uint380_t(x : std_logic_vector) return uint380_t;
subtype int380_t is signed(379 downto 0);
constant int380_t_SLV_LEN : integer := 380;
function int380_t_to_slv(x : int380_t) return std_logic_vector;
function slv_to_int380_t(x : std_logic_vector) return int380_t;
subtype uint381_t is unsigned(380 downto 0);
constant uint381_t_SLV_LEN : integer := 381;
function uint381_t_to_slv(x : uint381_t) return std_logic_vector;
function slv_to_uint381_t(x : std_logic_vector) return uint381_t;
subtype int381_t is signed(380 downto 0);
constant int381_t_SLV_LEN : integer := 381;
function int381_t_to_slv(x : int381_t) return std_logic_vector;
function slv_to_int381_t(x : std_logic_vector) return int381_t;
subtype uint382_t is unsigned(381 downto 0);
constant uint382_t_SLV_LEN : integer := 382;
function uint382_t_to_slv(x : uint382_t) return std_logic_vector;
function slv_to_uint382_t(x : std_logic_vector) return uint382_t;
subtype int382_t is signed(381 downto 0);
constant int382_t_SLV_LEN : integer := 382;
function int382_t_to_slv(x : int382_t) return std_logic_vector;
function slv_to_int382_t(x : std_logic_vector) return int382_t;
subtype uint383_t is unsigned(382 downto 0);
constant uint383_t_SLV_LEN : integer := 383;
function uint383_t_to_slv(x : uint383_t) return std_logic_vector;
function slv_to_uint383_t(x : std_logic_vector) return uint383_t;
subtype int383_t is signed(382 downto 0);
constant int383_t_SLV_LEN : integer := 383;
function int383_t_to_slv(x : int383_t) return std_logic_vector;
function slv_to_int383_t(x : std_logic_vector) return int383_t;
subtype uint384_t is unsigned(383 downto 0);
constant uint384_t_SLV_LEN : integer := 384;
function uint384_t_to_slv(x : uint384_t) return std_logic_vector;
function slv_to_uint384_t(x : std_logic_vector) return uint384_t;
subtype int384_t is signed(383 downto 0);
constant int384_t_SLV_LEN : integer := 384;
function int384_t_to_slv(x : int384_t) return std_logic_vector;
function slv_to_int384_t(x : std_logic_vector) return int384_t;
subtype uint385_t is unsigned(384 downto 0);
constant uint385_t_SLV_LEN : integer := 385;
function uint385_t_to_slv(x : uint385_t) return std_logic_vector;
function slv_to_uint385_t(x : std_logic_vector) return uint385_t;
subtype int385_t is signed(384 downto 0);
constant int385_t_SLV_LEN : integer := 385;
function int385_t_to_slv(x : int385_t) return std_logic_vector;
function slv_to_int385_t(x : std_logic_vector) return int385_t;
subtype uint386_t is unsigned(385 downto 0);
constant uint386_t_SLV_LEN : integer := 386;
function uint386_t_to_slv(x : uint386_t) return std_logic_vector;
function slv_to_uint386_t(x : std_logic_vector) return uint386_t;
subtype int386_t is signed(385 downto 0);
constant int386_t_SLV_LEN : integer := 386;
function int386_t_to_slv(x : int386_t) return std_logic_vector;
function slv_to_int386_t(x : std_logic_vector) return int386_t;
subtype uint387_t is unsigned(386 downto 0);
constant uint387_t_SLV_LEN : integer := 387;
function uint387_t_to_slv(x : uint387_t) return std_logic_vector;
function slv_to_uint387_t(x : std_logic_vector) return uint387_t;
subtype int387_t is signed(386 downto 0);
constant int387_t_SLV_LEN : integer := 387;
function int387_t_to_slv(x : int387_t) return std_logic_vector;
function slv_to_int387_t(x : std_logic_vector) return int387_t;
subtype uint388_t is unsigned(387 downto 0);
constant uint388_t_SLV_LEN : integer := 388;
function uint388_t_to_slv(x : uint388_t) return std_logic_vector;
function slv_to_uint388_t(x : std_logic_vector) return uint388_t;
subtype int388_t is signed(387 downto 0);
constant int388_t_SLV_LEN : integer := 388;
function int388_t_to_slv(x : int388_t) return std_logic_vector;
function slv_to_int388_t(x : std_logic_vector) return int388_t;
subtype uint389_t is unsigned(388 downto 0);
constant uint389_t_SLV_LEN : integer := 389;
function uint389_t_to_slv(x : uint389_t) return std_logic_vector;
function slv_to_uint389_t(x : std_logic_vector) return uint389_t;
subtype int389_t is signed(388 downto 0);
constant int389_t_SLV_LEN : integer := 389;
function int389_t_to_slv(x : int389_t) return std_logic_vector;
function slv_to_int389_t(x : std_logic_vector) return int389_t;
subtype uint390_t is unsigned(389 downto 0);
constant uint390_t_SLV_LEN : integer := 390;
function uint390_t_to_slv(x : uint390_t) return std_logic_vector;
function slv_to_uint390_t(x : std_logic_vector) return uint390_t;
subtype int390_t is signed(389 downto 0);
constant int390_t_SLV_LEN : integer := 390;
function int390_t_to_slv(x : int390_t) return std_logic_vector;
function slv_to_int390_t(x : std_logic_vector) return int390_t;
subtype uint391_t is unsigned(390 downto 0);
constant uint391_t_SLV_LEN : integer := 391;
function uint391_t_to_slv(x : uint391_t) return std_logic_vector;
function slv_to_uint391_t(x : std_logic_vector) return uint391_t;
subtype int391_t is signed(390 downto 0);
constant int391_t_SLV_LEN : integer := 391;
function int391_t_to_slv(x : int391_t) return std_logic_vector;
function slv_to_int391_t(x : std_logic_vector) return int391_t;
subtype uint392_t is unsigned(391 downto 0);
constant uint392_t_SLV_LEN : integer := 392;
function uint392_t_to_slv(x : uint392_t) return std_logic_vector;
function slv_to_uint392_t(x : std_logic_vector) return uint392_t;
subtype int392_t is signed(391 downto 0);
constant int392_t_SLV_LEN : integer := 392;
function int392_t_to_slv(x : int392_t) return std_logic_vector;
function slv_to_int392_t(x : std_logic_vector) return int392_t;
subtype uint393_t is unsigned(392 downto 0);
constant uint393_t_SLV_LEN : integer := 393;
function uint393_t_to_slv(x : uint393_t) return std_logic_vector;
function slv_to_uint393_t(x : std_logic_vector) return uint393_t;
subtype int393_t is signed(392 downto 0);
constant int393_t_SLV_LEN : integer := 393;
function int393_t_to_slv(x : int393_t) return std_logic_vector;
function slv_to_int393_t(x : std_logic_vector) return int393_t;
subtype uint394_t is unsigned(393 downto 0);
constant uint394_t_SLV_LEN : integer := 394;
function uint394_t_to_slv(x : uint394_t) return std_logic_vector;
function slv_to_uint394_t(x : std_logic_vector) return uint394_t;
subtype int394_t is signed(393 downto 0);
constant int394_t_SLV_LEN : integer := 394;
function int394_t_to_slv(x : int394_t) return std_logic_vector;
function slv_to_int394_t(x : std_logic_vector) return int394_t;
subtype uint395_t is unsigned(394 downto 0);
constant uint395_t_SLV_LEN : integer := 395;
function uint395_t_to_slv(x : uint395_t) return std_logic_vector;
function slv_to_uint395_t(x : std_logic_vector) return uint395_t;
subtype int395_t is signed(394 downto 0);
constant int395_t_SLV_LEN : integer := 395;
function int395_t_to_slv(x : int395_t) return std_logic_vector;
function slv_to_int395_t(x : std_logic_vector) return int395_t;
subtype uint396_t is unsigned(395 downto 0);
constant uint396_t_SLV_LEN : integer := 396;
function uint396_t_to_slv(x : uint396_t) return std_logic_vector;
function slv_to_uint396_t(x : std_logic_vector) return uint396_t;
subtype int396_t is signed(395 downto 0);
constant int396_t_SLV_LEN : integer := 396;
function int396_t_to_slv(x : int396_t) return std_logic_vector;
function slv_to_int396_t(x : std_logic_vector) return int396_t;
subtype uint397_t is unsigned(396 downto 0);
constant uint397_t_SLV_LEN : integer := 397;
function uint397_t_to_slv(x : uint397_t) return std_logic_vector;
function slv_to_uint397_t(x : std_logic_vector) return uint397_t;
subtype int397_t is signed(396 downto 0);
constant int397_t_SLV_LEN : integer := 397;
function int397_t_to_slv(x : int397_t) return std_logic_vector;
function slv_to_int397_t(x : std_logic_vector) return int397_t;
subtype uint398_t is unsigned(397 downto 0);
constant uint398_t_SLV_LEN : integer := 398;
function uint398_t_to_slv(x : uint398_t) return std_logic_vector;
function slv_to_uint398_t(x : std_logic_vector) return uint398_t;
subtype int398_t is signed(397 downto 0);
constant int398_t_SLV_LEN : integer := 398;
function int398_t_to_slv(x : int398_t) return std_logic_vector;
function slv_to_int398_t(x : std_logic_vector) return int398_t;
subtype uint399_t is unsigned(398 downto 0);
constant uint399_t_SLV_LEN : integer := 399;
function uint399_t_to_slv(x : uint399_t) return std_logic_vector;
function slv_to_uint399_t(x : std_logic_vector) return uint399_t;
subtype int399_t is signed(398 downto 0);
constant int399_t_SLV_LEN : integer := 399;
function int399_t_to_slv(x : int399_t) return std_logic_vector;
function slv_to_int399_t(x : std_logic_vector) return int399_t;
subtype uint400_t is unsigned(399 downto 0);
constant uint400_t_SLV_LEN : integer := 400;
function uint400_t_to_slv(x : uint400_t) return std_logic_vector;
function slv_to_uint400_t(x : std_logic_vector) return uint400_t;
subtype int400_t is signed(399 downto 0);
constant int400_t_SLV_LEN : integer := 400;
function int400_t_to_slv(x : int400_t) return std_logic_vector;
function slv_to_int400_t(x : std_logic_vector) return int400_t;
subtype uint401_t is unsigned(400 downto 0);
constant uint401_t_SLV_LEN : integer := 401;
function uint401_t_to_slv(x : uint401_t) return std_logic_vector;
function slv_to_uint401_t(x : std_logic_vector) return uint401_t;
subtype int401_t is signed(400 downto 0);
constant int401_t_SLV_LEN : integer := 401;
function int401_t_to_slv(x : int401_t) return std_logic_vector;
function slv_to_int401_t(x : std_logic_vector) return int401_t;
subtype uint402_t is unsigned(401 downto 0);
constant uint402_t_SLV_LEN : integer := 402;
function uint402_t_to_slv(x : uint402_t) return std_logic_vector;
function slv_to_uint402_t(x : std_logic_vector) return uint402_t;
subtype int402_t is signed(401 downto 0);
constant int402_t_SLV_LEN : integer := 402;
function int402_t_to_slv(x : int402_t) return std_logic_vector;
function slv_to_int402_t(x : std_logic_vector) return int402_t;
subtype uint403_t is unsigned(402 downto 0);
constant uint403_t_SLV_LEN : integer := 403;
function uint403_t_to_slv(x : uint403_t) return std_logic_vector;
function slv_to_uint403_t(x : std_logic_vector) return uint403_t;
subtype int403_t is signed(402 downto 0);
constant int403_t_SLV_LEN : integer := 403;
function int403_t_to_slv(x : int403_t) return std_logic_vector;
function slv_to_int403_t(x : std_logic_vector) return int403_t;
subtype uint404_t is unsigned(403 downto 0);
constant uint404_t_SLV_LEN : integer := 404;
function uint404_t_to_slv(x : uint404_t) return std_logic_vector;
function slv_to_uint404_t(x : std_logic_vector) return uint404_t;
subtype int404_t is signed(403 downto 0);
constant int404_t_SLV_LEN : integer := 404;
function int404_t_to_slv(x : int404_t) return std_logic_vector;
function slv_to_int404_t(x : std_logic_vector) return int404_t;
subtype uint405_t is unsigned(404 downto 0);
constant uint405_t_SLV_LEN : integer := 405;
function uint405_t_to_slv(x : uint405_t) return std_logic_vector;
function slv_to_uint405_t(x : std_logic_vector) return uint405_t;
subtype int405_t is signed(404 downto 0);
constant int405_t_SLV_LEN : integer := 405;
function int405_t_to_slv(x : int405_t) return std_logic_vector;
function slv_to_int405_t(x : std_logic_vector) return int405_t;
subtype uint406_t is unsigned(405 downto 0);
constant uint406_t_SLV_LEN : integer := 406;
function uint406_t_to_slv(x : uint406_t) return std_logic_vector;
function slv_to_uint406_t(x : std_logic_vector) return uint406_t;
subtype int406_t is signed(405 downto 0);
constant int406_t_SLV_LEN : integer := 406;
function int406_t_to_slv(x : int406_t) return std_logic_vector;
function slv_to_int406_t(x : std_logic_vector) return int406_t;
subtype uint407_t is unsigned(406 downto 0);
constant uint407_t_SLV_LEN : integer := 407;
function uint407_t_to_slv(x : uint407_t) return std_logic_vector;
function slv_to_uint407_t(x : std_logic_vector) return uint407_t;
subtype int407_t is signed(406 downto 0);
constant int407_t_SLV_LEN : integer := 407;
function int407_t_to_slv(x : int407_t) return std_logic_vector;
function slv_to_int407_t(x : std_logic_vector) return int407_t;
subtype uint408_t is unsigned(407 downto 0);
constant uint408_t_SLV_LEN : integer := 408;
function uint408_t_to_slv(x : uint408_t) return std_logic_vector;
function slv_to_uint408_t(x : std_logic_vector) return uint408_t;
subtype int408_t is signed(407 downto 0);
constant int408_t_SLV_LEN : integer := 408;
function int408_t_to_slv(x : int408_t) return std_logic_vector;
function slv_to_int408_t(x : std_logic_vector) return int408_t;
subtype uint409_t is unsigned(408 downto 0);
constant uint409_t_SLV_LEN : integer := 409;
function uint409_t_to_slv(x : uint409_t) return std_logic_vector;
function slv_to_uint409_t(x : std_logic_vector) return uint409_t;
subtype int409_t is signed(408 downto 0);
constant int409_t_SLV_LEN : integer := 409;
function int409_t_to_slv(x : int409_t) return std_logic_vector;
function slv_to_int409_t(x : std_logic_vector) return int409_t;
subtype uint410_t is unsigned(409 downto 0);
constant uint410_t_SLV_LEN : integer := 410;
function uint410_t_to_slv(x : uint410_t) return std_logic_vector;
function slv_to_uint410_t(x : std_logic_vector) return uint410_t;
subtype int410_t is signed(409 downto 0);
constant int410_t_SLV_LEN : integer := 410;
function int410_t_to_slv(x : int410_t) return std_logic_vector;
function slv_to_int410_t(x : std_logic_vector) return int410_t;
subtype uint411_t is unsigned(410 downto 0);
constant uint411_t_SLV_LEN : integer := 411;
function uint411_t_to_slv(x : uint411_t) return std_logic_vector;
function slv_to_uint411_t(x : std_logic_vector) return uint411_t;
subtype int411_t is signed(410 downto 0);
constant int411_t_SLV_LEN : integer := 411;
function int411_t_to_slv(x : int411_t) return std_logic_vector;
function slv_to_int411_t(x : std_logic_vector) return int411_t;
subtype uint412_t is unsigned(411 downto 0);
constant uint412_t_SLV_LEN : integer := 412;
function uint412_t_to_slv(x : uint412_t) return std_logic_vector;
function slv_to_uint412_t(x : std_logic_vector) return uint412_t;
subtype int412_t is signed(411 downto 0);
constant int412_t_SLV_LEN : integer := 412;
function int412_t_to_slv(x : int412_t) return std_logic_vector;
function slv_to_int412_t(x : std_logic_vector) return int412_t;
subtype uint413_t is unsigned(412 downto 0);
constant uint413_t_SLV_LEN : integer := 413;
function uint413_t_to_slv(x : uint413_t) return std_logic_vector;
function slv_to_uint413_t(x : std_logic_vector) return uint413_t;
subtype int413_t is signed(412 downto 0);
constant int413_t_SLV_LEN : integer := 413;
function int413_t_to_slv(x : int413_t) return std_logic_vector;
function slv_to_int413_t(x : std_logic_vector) return int413_t;
subtype uint414_t is unsigned(413 downto 0);
constant uint414_t_SLV_LEN : integer := 414;
function uint414_t_to_slv(x : uint414_t) return std_logic_vector;
function slv_to_uint414_t(x : std_logic_vector) return uint414_t;
subtype int414_t is signed(413 downto 0);
constant int414_t_SLV_LEN : integer := 414;
function int414_t_to_slv(x : int414_t) return std_logic_vector;
function slv_to_int414_t(x : std_logic_vector) return int414_t;
subtype uint415_t is unsigned(414 downto 0);
constant uint415_t_SLV_LEN : integer := 415;
function uint415_t_to_slv(x : uint415_t) return std_logic_vector;
function slv_to_uint415_t(x : std_logic_vector) return uint415_t;
subtype int415_t is signed(414 downto 0);
constant int415_t_SLV_LEN : integer := 415;
function int415_t_to_slv(x : int415_t) return std_logic_vector;
function slv_to_int415_t(x : std_logic_vector) return int415_t;
subtype uint416_t is unsigned(415 downto 0);
constant uint416_t_SLV_LEN : integer := 416;
function uint416_t_to_slv(x : uint416_t) return std_logic_vector;
function slv_to_uint416_t(x : std_logic_vector) return uint416_t;
subtype int416_t is signed(415 downto 0);
constant int416_t_SLV_LEN : integer := 416;
function int416_t_to_slv(x : int416_t) return std_logic_vector;
function slv_to_int416_t(x : std_logic_vector) return int416_t;
subtype uint417_t is unsigned(416 downto 0);
constant uint417_t_SLV_LEN : integer := 417;
function uint417_t_to_slv(x : uint417_t) return std_logic_vector;
function slv_to_uint417_t(x : std_logic_vector) return uint417_t;
subtype int417_t is signed(416 downto 0);
constant int417_t_SLV_LEN : integer := 417;
function int417_t_to_slv(x : int417_t) return std_logic_vector;
function slv_to_int417_t(x : std_logic_vector) return int417_t;
subtype uint418_t is unsigned(417 downto 0);
constant uint418_t_SLV_LEN : integer := 418;
function uint418_t_to_slv(x : uint418_t) return std_logic_vector;
function slv_to_uint418_t(x : std_logic_vector) return uint418_t;
subtype int418_t is signed(417 downto 0);
constant int418_t_SLV_LEN : integer := 418;
function int418_t_to_slv(x : int418_t) return std_logic_vector;
function slv_to_int418_t(x : std_logic_vector) return int418_t;
subtype uint419_t is unsigned(418 downto 0);
constant uint419_t_SLV_LEN : integer := 419;
function uint419_t_to_slv(x : uint419_t) return std_logic_vector;
function slv_to_uint419_t(x : std_logic_vector) return uint419_t;
subtype int419_t is signed(418 downto 0);
constant int419_t_SLV_LEN : integer := 419;
function int419_t_to_slv(x : int419_t) return std_logic_vector;
function slv_to_int419_t(x : std_logic_vector) return int419_t;
subtype uint420_t is unsigned(419 downto 0);
constant uint420_t_SLV_LEN : integer := 420;
function uint420_t_to_slv(x : uint420_t) return std_logic_vector;
function slv_to_uint420_t(x : std_logic_vector) return uint420_t;
subtype int420_t is signed(419 downto 0);
constant int420_t_SLV_LEN : integer := 420;
function int420_t_to_slv(x : int420_t) return std_logic_vector;
function slv_to_int420_t(x : std_logic_vector) return int420_t;
subtype uint421_t is unsigned(420 downto 0);
constant uint421_t_SLV_LEN : integer := 421;
function uint421_t_to_slv(x : uint421_t) return std_logic_vector;
function slv_to_uint421_t(x : std_logic_vector) return uint421_t;
subtype int421_t is signed(420 downto 0);
constant int421_t_SLV_LEN : integer := 421;
function int421_t_to_slv(x : int421_t) return std_logic_vector;
function slv_to_int421_t(x : std_logic_vector) return int421_t;
subtype uint422_t is unsigned(421 downto 0);
constant uint422_t_SLV_LEN : integer := 422;
function uint422_t_to_slv(x : uint422_t) return std_logic_vector;
function slv_to_uint422_t(x : std_logic_vector) return uint422_t;
subtype int422_t is signed(421 downto 0);
constant int422_t_SLV_LEN : integer := 422;
function int422_t_to_slv(x : int422_t) return std_logic_vector;
function slv_to_int422_t(x : std_logic_vector) return int422_t;
subtype uint423_t is unsigned(422 downto 0);
constant uint423_t_SLV_LEN : integer := 423;
function uint423_t_to_slv(x : uint423_t) return std_logic_vector;
function slv_to_uint423_t(x : std_logic_vector) return uint423_t;
subtype int423_t is signed(422 downto 0);
constant int423_t_SLV_LEN : integer := 423;
function int423_t_to_slv(x : int423_t) return std_logic_vector;
function slv_to_int423_t(x : std_logic_vector) return int423_t;
subtype uint424_t is unsigned(423 downto 0);
constant uint424_t_SLV_LEN : integer := 424;
function uint424_t_to_slv(x : uint424_t) return std_logic_vector;
function slv_to_uint424_t(x : std_logic_vector) return uint424_t;
subtype int424_t is signed(423 downto 0);
constant int424_t_SLV_LEN : integer := 424;
function int424_t_to_slv(x : int424_t) return std_logic_vector;
function slv_to_int424_t(x : std_logic_vector) return int424_t;
subtype uint425_t is unsigned(424 downto 0);
constant uint425_t_SLV_LEN : integer := 425;
function uint425_t_to_slv(x : uint425_t) return std_logic_vector;
function slv_to_uint425_t(x : std_logic_vector) return uint425_t;
subtype int425_t is signed(424 downto 0);
constant int425_t_SLV_LEN : integer := 425;
function int425_t_to_slv(x : int425_t) return std_logic_vector;
function slv_to_int425_t(x : std_logic_vector) return int425_t;
subtype uint426_t is unsigned(425 downto 0);
constant uint426_t_SLV_LEN : integer := 426;
function uint426_t_to_slv(x : uint426_t) return std_logic_vector;
function slv_to_uint426_t(x : std_logic_vector) return uint426_t;
subtype int426_t is signed(425 downto 0);
constant int426_t_SLV_LEN : integer := 426;
function int426_t_to_slv(x : int426_t) return std_logic_vector;
function slv_to_int426_t(x : std_logic_vector) return int426_t;
subtype uint427_t is unsigned(426 downto 0);
constant uint427_t_SLV_LEN : integer := 427;
function uint427_t_to_slv(x : uint427_t) return std_logic_vector;
function slv_to_uint427_t(x : std_logic_vector) return uint427_t;
subtype int427_t is signed(426 downto 0);
constant int427_t_SLV_LEN : integer := 427;
function int427_t_to_slv(x : int427_t) return std_logic_vector;
function slv_to_int427_t(x : std_logic_vector) return int427_t;
subtype uint428_t is unsigned(427 downto 0);
constant uint428_t_SLV_LEN : integer := 428;
function uint428_t_to_slv(x : uint428_t) return std_logic_vector;
function slv_to_uint428_t(x : std_logic_vector) return uint428_t;
subtype int428_t is signed(427 downto 0);
constant int428_t_SLV_LEN : integer := 428;
function int428_t_to_slv(x : int428_t) return std_logic_vector;
function slv_to_int428_t(x : std_logic_vector) return int428_t;
subtype uint429_t is unsigned(428 downto 0);
constant uint429_t_SLV_LEN : integer := 429;
function uint429_t_to_slv(x : uint429_t) return std_logic_vector;
function slv_to_uint429_t(x : std_logic_vector) return uint429_t;
subtype int429_t is signed(428 downto 0);
constant int429_t_SLV_LEN : integer := 429;
function int429_t_to_slv(x : int429_t) return std_logic_vector;
function slv_to_int429_t(x : std_logic_vector) return int429_t;
subtype uint430_t is unsigned(429 downto 0);
constant uint430_t_SLV_LEN : integer := 430;
function uint430_t_to_slv(x : uint430_t) return std_logic_vector;
function slv_to_uint430_t(x : std_logic_vector) return uint430_t;
subtype int430_t is signed(429 downto 0);
constant int430_t_SLV_LEN : integer := 430;
function int430_t_to_slv(x : int430_t) return std_logic_vector;
function slv_to_int430_t(x : std_logic_vector) return int430_t;
subtype uint431_t is unsigned(430 downto 0);
constant uint431_t_SLV_LEN : integer := 431;
function uint431_t_to_slv(x : uint431_t) return std_logic_vector;
function slv_to_uint431_t(x : std_logic_vector) return uint431_t;
subtype int431_t is signed(430 downto 0);
constant int431_t_SLV_LEN : integer := 431;
function int431_t_to_slv(x : int431_t) return std_logic_vector;
function slv_to_int431_t(x : std_logic_vector) return int431_t;
subtype uint432_t is unsigned(431 downto 0);
constant uint432_t_SLV_LEN : integer := 432;
function uint432_t_to_slv(x : uint432_t) return std_logic_vector;
function slv_to_uint432_t(x : std_logic_vector) return uint432_t;
subtype int432_t is signed(431 downto 0);
constant int432_t_SLV_LEN : integer := 432;
function int432_t_to_slv(x : int432_t) return std_logic_vector;
function slv_to_int432_t(x : std_logic_vector) return int432_t;
subtype uint433_t is unsigned(432 downto 0);
constant uint433_t_SLV_LEN : integer := 433;
function uint433_t_to_slv(x : uint433_t) return std_logic_vector;
function slv_to_uint433_t(x : std_logic_vector) return uint433_t;
subtype int433_t is signed(432 downto 0);
constant int433_t_SLV_LEN : integer := 433;
function int433_t_to_slv(x : int433_t) return std_logic_vector;
function slv_to_int433_t(x : std_logic_vector) return int433_t;
subtype uint434_t is unsigned(433 downto 0);
constant uint434_t_SLV_LEN : integer := 434;
function uint434_t_to_slv(x : uint434_t) return std_logic_vector;
function slv_to_uint434_t(x : std_logic_vector) return uint434_t;
subtype int434_t is signed(433 downto 0);
constant int434_t_SLV_LEN : integer := 434;
function int434_t_to_slv(x : int434_t) return std_logic_vector;
function slv_to_int434_t(x : std_logic_vector) return int434_t;
subtype uint435_t is unsigned(434 downto 0);
constant uint435_t_SLV_LEN : integer := 435;
function uint435_t_to_slv(x : uint435_t) return std_logic_vector;
function slv_to_uint435_t(x : std_logic_vector) return uint435_t;
subtype int435_t is signed(434 downto 0);
constant int435_t_SLV_LEN : integer := 435;
function int435_t_to_slv(x : int435_t) return std_logic_vector;
function slv_to_int435_t(x : std_logic_vector) return int435_t;
subtype uint436_t is unsigned(435 downto 0);
constant uint436_t_SLV_LEN : integer := 436;
function uint436_t_to_slv(x : uint436_t) return std_logic_vector;
function slv_to_uint436_t(x : std_logic_vector) return uint436_t;
subtype int436_t is signed(435 downto 0);
constant int436_t_SLV_LEN : integer := 436;
function int436_t_to_slv(x : int436_t) return std_logic_vector;
function slv_to_int436_t(x : std_logic_vector) return int436_t;
subtype uint437_t is unsigned(436 downto 0);
constant uint437_t_SLV_LEN : integer := 437;
function uint437_t_to_slv(x : uint437_t) return std_logic_vector;
function slv_to_uint437_t(x : std_logic_vector) return uint437_t;
subtype int437_t is signed(436 downto 0);
constant int437_t_SLV_LEN : integer := 437;
function int437_t_to_slv(x : int437_t) return std_logic_vector;
function slv_to_int437_t(x : std_logic_vector) return int437_t;
subtype uint438_t is unsigned(437 downto 0);
constant uint438_t_SLV_LEN : integer := 438;
function uint438_t_to_slv(x : uint438_t) return std_logic_vector;
function slv_to_uint438_t(x : std_logic_vector) return uint438_t;
subtype int438_t is signed(437 downto 0);
constant int438_t_SLV_LEN : integer := 438;
function int438_t_to_slv(x : int438_t) return std_logic_vector;
function slv_to_int438_t(x : std_logic_vector) return int438_t;
subtype uint439_t is unsigned(438 downto 0);
constant uint439_t_SLV_LEN : integer := 439;
function uint439_t_to_slv(x : uint439_t) return std_logic_vector;
function slv_to_uint439_t(x : std_logic_vector) return uint439_t;
subtype int439_t is signed(438 downto 0);
constant int439_t_SLV_LEN : integer := 439;
function int439_t_to_slv(x : int439_t) return std_logic_vector;
function slv_to_int439_t(x : std_logic_vector) return int439_t;
subtype uint440_t is unsigned(439 downto 0);
constant uint440_t_SLV_LEN : integer := 440;
function uint440_t_to_slv(x : uint440_t) return std_logic_vector;
function slv_to_uint440_t(x : std_logic_vector) return uint440_t;
subtype int440_t is signed(439 downto 0);
constant int440_t_SLV_LEN : integer := 440;
function int440_t_to_slv(x : int440_t) return std_logic_vector;
function slv_to_int440_t(x : std_logic_vector) return int440_t;
subtype uint441_t is unsigned(440 downto 0);
constant uint441_t_SLV_LEN : integer := 441;
function uint441_t_to_slv(x : uint441_t) return std_logic_vector;
function slv_to_uint441_t(x : std_logic_vector) return uint441_t;
subtype int441_t is signed(440 downto 0);
constant int441_t_SLV_LEN : integer := 441;
function int441_t_to_slv(x : int441_t) return std_logic_vector;
function slv_to_int441_t(x : std_logic_vector) return int441_t;
subtype uint442_t is unsigned(441 downto 0);
constant uint442_t_SLV_LEN : integer := 442;
function uint442_t_to_slv(x : uint442_t) return std_logic_vector;
function slv_to_uint442_t(x : std_logic_vector) return uint442_t;
subtype int442_t is signed(441 downto 0);
constant int442_t_SLV_LEN : integer := 442;
function int442_t_to_slv(x : int442_t) return std_logic_vector;
function slv_to_int442_t(x : std_logic_vector) return int442_t;
subtype uint443_t is unsigned(442 downto 0);
constant uint443_t_SLV_LEN : integer := 443;
function uint443_t_to_slv(x : uint443_t) return std_logic_vector;
function slv_to_uint443_t(x : std_logic_vector) return uint443_t;
subtype int443_t is signed(442 downto 0);
constant int443_t_SLV_LEN : integer := 443;
function int443_t_to_slv(x : int443_t) return std_logic_vector;
function slv_to_int443_t(x : std_logic_vector) return int443_t;
subtype uint444_t is unsigned(443 downto 0);
constant uint444_t_SLV_LEN : integer := 444;
function uint444_t_to_slv(x : uint444_t) return std_logic_vector;
function slv_to_uint444_t(x : std_logic_vector) return uint444_t;
subtype int444_t is signed(443 downto 0);
constant int444_t_SLV_LEN : integer := 444;
function int444_t_to_slv(x : int444_t) return std_logic_vector;
function slv_to_int444_t(x : std_logic_vector) return int444_t;
subtype uint445_t is unsigned(444 downto 0);
constant uint445_t_SLV_LEN : integer := 445;
function uint445_t_to_slv(x : uint445_t) return std_logic_vector;
function slv_to_uint445_t(x : std_logic_vector) return uint445_t;
subtype int445_t is signed(444 downto 0);
constant int445_t_SLV_LEN : integer := 445;
function int445_t_to_slv(x : int445_t) return std_logic_vector;
function slv_to_int445_t(x : std_logic_vector) return int445_t;
subtype uint446_t is unsigned(445 downto 0);
constant uint446_t_SLV_LEN : integer := 446;
function uint446_t_to_slv(x : uint446_t) return std_logic_vector;
function slv_to_uint446_t(x : std_logic_vector) return uint446_t;
subtype int446_t is signed(445 downto 0);
constant int446_t_SLV_LEN : integer := 446;
function int446_t_to_slv(x : int446_t) return std_logic_vector;
function slv_to_int446_t(x : std_logic_vector) return int446_t;
subtype uint447_t is unsigned(446 downto 0);
constant uint447_t_SLV_LEN : integer := 447;
function uint447_t_to_slv(x : uint447_t) return std_logic_vector;
function slv_to_uint447_t(x : std_logic_vector) return uint447_t;
subtype int447_t is signed(446 downto 0);
constant int447_t_SLV_LEN : integer := 447;
function int447_t_to_slv(x : int447_t) return std_logic_vector;
function slv_to_int447_t(x : std_logic_vector) return int447_t;
subtype uint448_t is unsigned(447 downto 0);
constant uint448_t_SLV_LEN : integer := 448;
function uint448_t_to_slv(x : uint448_t) return std_logic_vector;
function slv_to_uint448_t(x : std_logic_vector) return uint448_t;
subtype int448_t is signed(447 downto 0);
constant int448_t_SLV_LEN : integer := 448;
function int448_t_to_slv(x : int448_t) return std_logic_vector;
function slv_to_int448_t(x : std_logic_vector) return int448_t;
subtype uint449_t is unsigned(448 downto 0);
constant uint449_t_SLV_LEN : integer := 449;
function uint449_t_to_slv(x : uint449_t) return std_logic_vector;
function slv_to_uint449_t(x : std_logic_vector) return uint449_t;
subtype int449_t is signed(448 downto 0);
constant int449_t_SLV_LEN : integer := 449;
function int449_t_to_slv(x : int449_t) return std_logic_vector;
function slv_to_int449_t(x : std_logic_vector) return int449_t;
subtype uint450_t is unsigned(449 downto 0);
constant uint450_t_SLV_LEN : integer := 450;
function uint450_t_to_slv(x : uint450_t) return std_logic_vector;
function slv_to_uint450_t(x : std_logic_vector) return uint450_t;
subtype int450_t is signed(449 downto 0);
constant int450_t_SLV_LEN : integer := 450;
function int450_t_to_slv(x : int450_t) return std_logic_vector;
function slv_to_int450_t(x : std_logic_vector) return int450_t;
subtype uint451_t is unsigned(450 downto 0);
constant uint451_t_SLV_LEN : integer := 451;
function uint451_t_to_slv(x : uint451_t) return std_logic_vector;
function slv_to_uint451_t(x : std_logic_vector) return uint451_t;
subtype int451_t is signed(450 downto 0);
constant int451_t_SLV_LEN : integer := 451;
function int451_t_to_slv(x : int451_t) return std_logic_vector;
function slv_to_int451_t(x : std_logic_vector) return int451_t;
subtype uint452_t is unsigned(451 downto 0);
constant uint452_t_SLV_LEN : integer := 452;
function uint452_t_to_slv(x : uint452_t) return std_logic_vector;
function slv_to_uint452_t(x : std_logic_vector) return uint452_t;
subtype int452_t is signed(451 downto 0);
constant int452_t_SLV_LEN : integer := 452;
function int452_t_to_slv(x : int452_t) return std_logic_vector;
function slv_to_int452_t(x : std_logic_vector) return int452_t;
subtype uint453_t is unsigned(452 downto 0);
constant uint453_t_SLV_LEN : integer := 453;
function uint453_t_to_slv(x : uint453_t) return std_logic_vector;
function slv_to_uint453_t(x : std_logic_vector) return uint453_t;
subtype int453_t is signed(452 downto 0);
constant int453_t_SLV_LEN : integer := 453;
function int453_t_to_slv(x : int453_t) return std_logic_vector;
function slv_to_int453_t(x : std_logic_vector) return int453_t;
subtype uint454_t is unsigned(453 downto 0);
constant uint454_t_SLV_LEN : integer := 454;
function uint454_t_to_slv(x : uint454_t) return std_logic_vector;
function slv_to_uint454_t(x : std_logic_vector) return uint454_t;
subtype int454_t is signed(453 downto 0);
constant int454_t_SLV_LEN : integer := 454;
function int454_t_to_slv(x : int454_t) return std_logic_vector;
function slv_to_int454_t(x : std_logic_vector) return int454_t;
subtype uint455_t is unsigned(454 downto 0);
constant uint455_t_SLV_LEN : integer := 455;
function uint455_t_to_slv(x : uint455_t) return std_logic_vector;
function slv_to_uint455_t(x : std_logic_vector) return uint455_t;
subtype int455_t is signed(454 downto 0);
constant int455_t_SLV_LEN : integer := 455;
function int455_t_to_slv(x : int455_t) return std_logic_vector;
function slv_to_int455_t(x : std_logic_vector) return int455_t;
subtype uint456_t is unsigned(455 downto 0);
constant uint456_t_SLV_LEN : integer := 456;
function uint456_t_to_slv(x : uint456_t) return std_logic_vector;
function slv_to_uint456_t(x : std_logic_vector) return uint456_t;
subtype int456_t is signed(455 downto 0);
constant int456_t_SLV_LEN : integer := 456;
function int456_t_to_slv(x : int456_t) return std_logic_vector;
function slv_to_int456_t(x : std_logic_vector) return int456_t;
subtype uint457_t is unsigned(456 downto 0);
constant uint457_t_SLV_LEN : integer := 457;
function uint457_t_to_slv(x : uint457_t) return std_logic_vector;
function slv_to_uint457_t(x : std_logic_vector) return uint457_t;
subtype int457_t is signed(456 downto 0);
constant int457_t_SLV_LEN : integer := 457;
function int457_t_to_slv(x : int457_t) return std_logic_vector;
function slv_to_int457_t(x : std_logic_vector) return int457_t;
subtype uint458_t is unsigned(457 downto 0);
constant uint458_t_SLV_LEN : integer := 458;
function uint458_t_to_slv(x : uint458_t) return std_logic_vector;
function slv_to_uint458_t(x : std_logic_vector) return uint458_t;
subtype int458_t is signed(457 downto 0);
constant int458_t_SLV_LEN : integer := 458;
function int458_t_to_slv(x : int458_t) return std_logic_vector;
function slv_to_int458_t(x : std_logic_vector) return int458_t;
subtype uint459_t is unsigned(458 downto 0);
constant uint459_t_SLV_LEN : integer := 459;
function uint459_t_to_slv(x : uint459_t) return std_logic_vector;
function slv_to_uint459_t(x : std_logic_vector) return uint459_t;
subtype int459_t is signed(458 downto 0);
constant int459_t_SLV_LEN : integer := 459;
function int459_t_to_slv(x : int459_t) return std_logic_vector;
function slv_to_int459_t(x : std_logic_vector) return int459_t;
subtype uint460_t is unsigned(459 downto 0);
constant uint460_t_SLV_LEN : integer := 460;
function uint460_t_to_slv(x : uint460_t) return std_logic_vector;
function slv_to_uint460_t(x : std_logic_vector) return uint460_t;
subtype int460_t is signed(459 downto 0);
constant int460_t_SLV_LEN : integer := 460;
function int460_t_to_slv(x : int460_t) return std_logic_vector;
function slv_to_int460_t(x : std_logic_vector) return int460_t;
subtype uint461_t is unsigned(460 downto 0);
constant uint461_t_SLV_LEN : integer := 461;
function uint461_t_to_slv(x : uint461_t) return std_logic_vector;
function slv_to_uint461_t(x : std_logic_vector) return uint461_t;
subtype int461_t is signed(460 downto 0);
constant int461_t_SLV_LEN : integer := 461;
function int461_t_to_slv(x : int461_t) return std_logic_vector;
function slv_to_int461_t(x : std_logic_vector) return int461_t;
subtype uint462_t is unsigned(461 downto 0);
constant uint462_t_SLV_LEN : integer := 462;
function uint462_t_to_slv(x : uint462_t) return std_logic_vector;
function slv_to_uint462_t(x : std_logic_vector) return uint462_t;
subtype int462_t is signed(461 downto 0);
constant int462_t_SLV_LEN : integer := 462;
function int462_t_to_slv(x : int462_t) return std_logic_vector;
function slv_to_int462_t(x : std_logic_vector) return int462_t;
subtype uint463_t is unsigned(462 downto 0);
constant uint463_t_SLV_LEN : integer := 463;
function uint463_t_to_slv(x : uint463_t) return std_logic_vector;
function slv_to_uint463_t(x : std_logic_vector) return uint463_t;
subtype int463_t is signed(462 downto 0);
constant int463_t_SLV_LEN : integer := 463;
function int463_t_to_slv(x : int463_t) return std_logic_vector;
function slv_to_int463_t(x : std_logic_vector) return int463_t;
subtype uint464_t is unsigned(463 downto 0);
constant uint464_t_SLV_LEN : integer := 464;
function uint464_t_to_slv(x : uint464_t) return std_logic_vector;
function slv_to_uint464_t(x : std_logic_vector) return uint464_t;
subtype int464_t is signed(463 downto 0);
constant int464_t_SLV_LEN : integer := 464;
function int464_t_to_slv(x : int464_t) return std_logic_vector;
function slv_to_int464_t(x : std_logic_vector) return int464_t;
subtype uint465_t is unsigned(464 downto 0);
constant uint465_t_SLV_LEN : integer := 465;
function uint465_t_to_slv(x : uint465_t) return std_logic_vector;
function slv_to_uint465_t(x : std_logic_vector) return uint465_t;
subtype int465_t is signed(464 downto 0);
constant int465_t_SLV_LEN : integer := 465;
function int465_t_to_slv(x : int465_t) return std_logic_vector;
function slv_to_int465_t(x : std_logic_vector) return int465_t;
subtype uint466_t is unsigned(465 downto 0);
constant uint466_t_SLV_LEN : integer := 466;
function uint466_t_to_slv(x : uint466_t) return std_logic_vector;
function slv_to_uint466_t(x : std_logic_vector) return uint466_t;
subtype int466_t is signed(465 downto 0);
constant int466_t_SLV_LEN : integer := 466;
function int466_t_to_slv(x : int466_t) return std_logic_vector;
function slv_to_int466_t(x : std_logic_vector) return int466_t;
subtype uint467_t is unsigned(466 downto 0);
constant uint467_t_SLV_LEN : integer := 467;
function uint467_t_to_slv(x : uint467_t) return std_logic_vector;
function slv_to_uint467_t(x : std_logic_vector) return uint467_t;
subtype int467_t is signed(466 downto 0);
constant int467_t_SLV_LEN : integer := 467;
function int467_t_to_slv(x : int467_t) return std_logic_vector;
function slv_to_int467_t(x : std_logic_vector) return int467_t;
subtype uint468_t is unsigned(467 downto 0);
constant uint468_t_SLV_LEN : integer := 468;
function uint468_t_to_slv(x : uint468_t) return std_logic_vector;
function slv_to_uint468_t(x : std_logic_vector) return uint468_t;
subtype int468_t is signed(467 downto 0);
constant int468_t_SLV_LEN : integer := 468;
function int468_t_to_slv(x : int468_t) return std_logic_vector;
function slv_to_int468_t(x : std_logic_vector) return int468_t;
subtype uint469_t is unsigned(468 downto 0);
constant uint469_t_SLV_LEN : integer := 469;
function uint469_t_to_slv(x : uint469_t) return std_logic_vector;
function slv_to_uint469_t(x : std_logic_vector) return uint469_t;
subtype int469_t is signed(468 downto 0);
constant int469_t_SLV_LEN : integer := 469;
function int469_t_to_slv(x : int469_t) return std_logic_vector;
function slv_to_int469_t(x : std_logic_vector) return int469_t;
subtype uint470_t is unsigned(469 downto 0);
constant uint470_t_SLV_LEN : integer := 470;
function uint470_t_to_slv(x : uint470_t) return std_logic_vector;
function slv_to_uint470_t(x : std_logic_vector) return uint470_t;
subtype int470_t is signed(469 downto 0);
constant int470_t_SLV_LEN : integer := 470;
function int470_t_to_slv(x : int470_t) return std_logic_vector;
function slv_to_int470_t(x : std_logic_vector) return int470_t;
subtype uint471_t is unsigned(470 downto 0);
constant uint471_t_SLV_LEN : integer := 471;
function uint471_t_to_slv(x : uint471_t) return std_logic_vector;
function slv_to_uint471_t(x : std_logic_vector) return uint471_t;
subtype int471_t is signed(470 downto 0);
constant int471_t_SLV_LEN : integer := 471;
function int471_t_to_slv(x : int471_t) return std_logic_vector;
function slv_to_int471_t(x : std_logic_vector) return int471_t;
subtype uint472_t is unsigned(471 downto 0);
constant uint472_t_SLV_LEN : integer := 472;
function uint472_t_to_slv(x : uint472_t) return std_logic_vector;
function slv_to_uint472_t(x : std_logic_vector) return uint472_t;
subtype int472_t is signed(471 downto 0);
constant int472_t_SLV_LEN : integer := 472;
function int472_t_to_slv(x : int472_t) return std_logic_vector;
function slv_to_int472_t(x : std_logic_vector) return int472_t;
subtype uint473_t is unsigned(472 downto 0);
constant uint473_t_SLV_LEN : integer := 473;
function uint473_t_to_slv(x : uint473_t) return std_logic_vector;
function slv_to_uint473_t(x : std_logic_vector) return uint473_t;
subtype int473_t is signed(472 downto 0);
constant int473_t_SLV_LEN : integer := 473;
function int473_t_to_slv(x : int473_t) return std_logic_vector;
function slv_to_int473_t(x : std_logic_vector) return int473_t;
subtype uint474_t is unsigned(473 downto 0);
constant uint474_t_SLV_LEN : integer := 474;
function uint474_t_to_slv(x : uint474_t) return std_logic_vector;
function slv_to_uint474_t(x : std_logic_vector) return uint474_t;
subtype int474_t is signed(473 downto 0);
constant int474_t_SLV_LEN : integer := 474;
function int474_t_to_slv(x : int474_t) return std_logic_vector;
function slv_to_int474_t(x : std_logic_vector) return int474_t;
subtype uint475_t is unsigned(474 downto 0);
constant uint475_t_SLV_LEN : integer := 475;
function uint475_t_to_slv(x : uint475_t) return std_logic_vector;
function slv_to_uint475_t(x : std_logic_vector) return uint475_t;
subtype int475_t is signed(474 downto 0);
constant int475_t_SLV_LEN : integer := 475;
function int475_t_to_slv(x : int475_t) return std_logic_vector;
function slv_to_int475_t(x : std_logic_vector) return int475_t;
subtype uint476_t is unsigned(475 downto 0);
constant uint476_t_SLV_LEN : integer := 476;
function uint476_t_to_slv(x : uint476_t) return std_logic_vector;
function slv_to_uint476_t(x : std_logic_vector) return uint476_t;
subtype int476_t is signed(475 downto 0);
constant int476_t_SLV_LEN : integer := 476;
function int476_t_to_slv(x : int476_t) return std_logic_vector;
function slv_to_int476_t(x : std_logic_vector) return int476_t;
subtype uint477_t is unsigned(476 downto 0);
constant uint477_t_SLV_LEN : integer := 477;
function uint477_t_to_slv(x : uint477_t) return std_logic_vector;
function slv_to_uint477_t(x : std_logic_vector) return uint477_t;
subtype int477_t is signed(476 downto 0);
constant int477_t_SLV_LEN : integer := 477;
function int477_t_to_slv(x : int477_t) return std_logic_vector;
function slv_to_int477_t(x : std_logic_vector) return int477_t;
subtype uint478_t is unsigned(477 downto 0);
constant uint478_t_SLV_LEN : integer := 478;
function uint478_t_to_slv(x : uint478_t) return std_logic_vector;
function slv_to_uint478_t(x : std_logic_vector) return uint478_t;
subtype int478_t is signed(477 downto 0);
constant int478_t_SLV_LEN : integer := 478;
function int478_t_to_slv(x : int478_t) return std_logic_vector;
function slv_to_int478_t(x : std_logic_vector) return int478_t;
subtype uint479_t is unsigned(478 downto 0);
constant uint479_t_SLV_LEN : integer := 479;
function uint479_t_to_slv(x : uint479_t) return std_logic_vector;
function slv_to_uint479_t(x : std_logic_vector) return uint479_t;
subtype int479_t is signed(478 downto 0);
constant int479_t_SLV_LEN : integer := 479;
function int479_t_to_slv(x : int479_t) return std_logic_vector;
function slv_to_int479_t(x : std_logic_vector) return int479_t;
subtype uint480_t is unsigned(479 downto 0);
constant uint480_t_SLV_LEN : integer := 480;
function uint480_t_to_slv(x : uint480_t) return std_logic_vector;
function slv_to_uint480_t(x : std_logic_vector) return uint480_t;
subtype int480_t is signed(479 downto 0);
constant int480_t_SLV_LEN : integer := 480;
function int480_t_to_slv(x : int480_t) return std_logic_vector;
function slv_to_int480_t(x : std_logic_vector) return int480_t;
subtype uint481_t is unsigned(480 downto 0);
constant uint481_t_SLV_LEN : integer := 481;
function uint481_t_to_slv(x : uint481_t) return std_logic_vector;
function slv_to_uint481_t(x : std_logic_vector) return uint481_t;
subtype int481_t is signed(480 downto 0);
constant int481_t_SLV_LEN : integer := 481;
function int481_t_to_slv(x : int481_t) return std_logic_vector;
function slv_to_int481_t(x : std_logic_vector) return int481_t;
subtype uint482_t is unsigned(481 downto 0);
constant uint482_t_SLV_LEN : integer := 482;
function uint482_t_to_slv(x : uint482_t) return std_logic_vector;
function slv_to_uint482_t(x : std_logic_vector) return uint482_t;
subtype int482_t is signed(481 downto 0);
constant int482_t_SLV_LEN : integer := 482;
function int482_t_to_slv(x : int482_t) return std_logic_vector;
function slv_to_int482_t(x : std_logic_vector) return int482_t;
subtype uint483_t is unsigned(482 downto 0);
constant uint483_t_SLV_LEN : integer := 483;
function uint483_t_to_slv(x : uint483_t) return std_logic_vector;
function slv_to_uint483_t(x : std_logic_vector) return uint483_t;
subtype int483_t is signed(482 downto 0);
constant int483_t_SLV_LEN : integer := 483;
function int483_t_to_slv(x : int483_t) return std_logic_vector;
function slv_to_int483_t(x : std_logic_vector) return int483_t;
subtype uint484_t is unsigned(483 downto 0);
constant uint484_t_SLV_LEN : integer := 484;
function uint484_t_to_slv(x : uint484_t) return std_logic_vector;
function slv_to_uint484_t(x : std_logic_vector) return uint484_t;
subtype int484_t is signed(483 downto 0);
constant int484_t_SLV_LEN : integer := 484;
function int484_t_to_slv(x : int484_t) return std_logic_vector;
function slv_to_int484_t(x : std_logic_vector) return int484_t;
subtype uint485_t is unsigned(484 downto 0);
constant uint485_t_SLV_LEN : integer := 485;
function uint485_t_to_slv(x : uint485_t) return std_logic_vector;
function slv_to_uint485_t(x : std_logic_vector) return uint485_t;
subtype int485_t is signed(484 downto 0);
constant int485_t_SLV_LEN : integer := 485;
function int485_t_to_slv(x : int485_t) return std_logic_vector;
function slv_to_int485_t(x : std_logic_vector) return int485_t;
subtype uint486_t is unsigned(485 downto 0);
constant uint486_t_SLV_LEN : integer := 486;
function uint486_t_to_slv(x : uint486_t) return std_logic_vector;
function slv_to_uint486_t(x : std_logic_vector) return uint486_t;
subtype int486_t is signed(485 downto 0);
constant int486_t_SLV_LEN : integer := 486;
function int486_t_to_slv(x : int486_t) return std_logic_vector;
function slv_to_int486_t(x : std_logic_vector) return int486_t;
subtype uint487_t is unsigned(486 downto 0);
constant uint487_t_SLV_LEN : integer := 487;
function uint487_t_to_slv(x : uint487_t) return std_logic_vector;
function slv_to_uint487_t(x : std_logic_vector) return uint487_t;
subtype int487_t is signed(486 downto 0);
constant int487_t_SLV_LEN : integer := 487;
function int487_t_to_slv(x : int487_t) return std_logic_vector;
function slv_to_int487_t(x : std_logic_vector) return int487_t;
subtype uint488_t is unsigned(487 downto 0);
constant uint488_t_SLV_LEN : integer := 488;
function uint488_t_to_slv(x : uint488_t) return std_logic_vector;
function slv_to_uint488_t(x : std_logic_vector) return uint488_t;
subtype int488_t is signed(487 downto 0);
constant int488_t_SLV_LEN : integer := 488;
function int488_t_to_slv(x : int488_t) return std_logic_vector;
function slv_to_int488_t(x : std_logic_vector) return int488_t;
subtype uint489_t is unsigned(488 downto 0);
constant uint489_t_SLV_LEN : integer := 489;
function uint489_t_to_slv(x : uint489_t) return std_logic_vector;
function slv_to_uint489_t(x : std_logic_vector) return uint489_t;
subtype int489_t is signed(488 downto 0);
constant int489_t_SLV_LEN : integer := 489;
function int489_t_to_slv(x : int489_t) return std_logic_vector;
function slv_to_int489_t(x : std_logic_vector) return int489_t;
subtype uint490_t is unsigned(489 downto 0);
constant uint490_t_SLV_LEN : integer := 490;
function uint490_t_to_slv(x : uint490_t) return std_logic_vector;
function slv_to_uint490_t(x : std_logic_vector) return uint490_t;
subtype int490_t is signed(489 downto 0);
constant int490_t_SLV_LEN : integer := 490;
function int490_t_to_slv(x : int490_t) return std_logic_vector;
function slv_to_int490_t(x : std_logic_vector) return int490_t;
subtype uint491_t is unsigned(490 downto 0);
constant uint491_t_SLV_LEN : integer := 491;
function uint491_t_to_slv(x : uint491_t) return std_logic_vector;
function slv_to_uint491_t(x : std_logic_vector) return uint491_t;
subtype int491_t is signed(490 downto 0);
constant int491_t_SLV_LEN : integer := 491;
function int491_t_to_slv(x : int491_t) return std_logic_vector;
function slv_to_int491_t(x : std_logic_vector) return int491_t;
subtype uint492_t is unsigned(491 downto 0);
constant uint492_t_SLV_LEN : integer := 492;
function uint492_t_to_slv(x : uint492_t) return std_logic_vector;
function slv_to_uint492_t(x : std_logic_vector) return uint492_t;
subtype int492_t is signed(491 downto 0);
constant int492_t_SLV_LEN : integer := 492;
function int492_t_to_slv(x : int492_t) return std_logic_vector;
function slv_to_int492_t(x : std_logic_vector) return int492_t;
subtype uint493_t is unsigned(492 downto 0);
constant uint493_t_SLV_LEN : integer := 493;
function uint493_t_to_slv(x : uint493_t) return std_logic_vector;
function slv_to_uint493_t(x : std_logic_vector) return uint493_t;
subtype int493_t is signed(492 downto 0);
constant int493_t_SLV_LEN : integer := 493;
function int493_t_to_slv(x : int493_t) return std_logic_vector;
function slv_to_int493_t(x : std_logic_vector) return int493_t;
subtype uint494_t is unsigned(493 downto 0);
constant uint494_t_SLV_LEN : integer := 494;
function uint494_t_to_slv(x : uint494_t) return std_logic_vector;
function slv_to_uint494_t(x : std_logic_vector) return uint494_t;
subtype int494_t is signed(493 downto 0);
constant int494_t_SLV_LEN : integer := 494;
function int494_t_to_slv(x : int494_t) return std_logic_vector;
function slv_to_int494_t(x : std_logic_vector) return int494_t;
subtype uint495_t is unsigned(494 downto 0);
constant uint495_t_SLV_LEN : integer := 495;
function uint495_t_to_slv(x : uint495_t) return std_logic_vector;
function slv_to_uint495_t(x : std_logic_vector) return uint495_t;
subtype int495_t is signed(494 downto 0);
constant int495_t_SLV_LEN : integer := 495;
function int495_t_to_slv(x : int495_t) return std_logic_vector;
function slv_to_int495_t(x : std_logic_vector) return int495_t;
subtype uint496_t is unsigned(495 downto 0);
constant uint496_t_SLV_LEN : integer := 496;
function uint496_t_to_slv(x : uint496_t) return std_logic_vector;
function slv_to_uint496_t(x : std_logic_vector) return uint496_t;
subtype int496_t is signed(495 downto 0);
constant int496_t_SLV_LEN : integer := 496;
function int496_t_to_slv(x : int496_t) return std_logic_vector;
function slv_to_int496_t(x : std_logic_vector) return int496_t;
subtype uint497_t is unsigned(496 downto 0);
constant uint497_t_SLV_LEN : integer := 497;
function uint497_t_to_slv(x : uint497_t) return std_logic_vector;
function slv_to_uint497_t(x : std_logic_vector) return uint497_t;
subtype int497_t is signed(496 downto 0);
constant int497_t_SLV_LEN : integer := 497;
function int497_t_to_slv(x : int497_t) return std_logic_vector;
function slv_to_int497_t(x : std_logic_vector) return int497_t;
subtype uint498_t is unsigned(497 downto 0);
constant uint498_t_SLV_LEN : integer := 498;
function uint498_t_to_slv(x : uint498_t) return std_logic_vector;
function slv_to_uint498_t(x : std_logic_vector) return uint498_t;
subtype int498_t is signed(497 downto 0);
constant int498_t_SLV_LEN : integer := 498;
function int498_t_to_slv(x : int498_t) return std_logic_vector;
function slv_to_int498_t(x : std_logic_vector) return int498_t;
subtype uint499_t is unsigned(498 downto 0);
constant uint499_t_SLV_LEN : integer := 499;
function uint499_t_to_slv(x : uint499_t) return std_logic_vector;
function slv_to_uint499_t(x : std_logic_vector) return uint499_t;
subtype int499_t is signed(498 downto 0);
constant int499_t_SLV_LEN : integer := 499;
function int499_t_to_slv(x : int499_t) return std_logic_vector;
function slv_to_int499_t(x : std_logic_vector) return int499_t;
subtype uint500_t is unsigned(499 downto 0);
constant uint500_t_SLV_LEN : integer := 500;
function uint500_t_to_slv(x : uint500_t) return std_logic_vector;
function slv_to_uint500_t(x : std_logic_vector) return uint500_t;
subtype int500_t is signed(499 downto 0);
constant int500_t_SLV_LEN : integer := 500;
function int500_t_to_slv(x : int500_t) return std_logic_vector;
function slv_to_int500_t(x : std_logic_vector) return int500_t;
subtype uint501_t is unsigned(500 downto 0);
constant uint501_t_SLV_LEN : integer := 501;
function uint501_t_to_slv(x : uint501_t) return std_logic_vector;
function slv_to_uint501_t(x : std_logic_vector) return uint501_t;
subtype int501_t is signed(500 downto 0);
constant int501_t_SLV_LEN : integer := 501;
function int501_t_to_slv(x : int501_t) return std_logic_vector;
function slv_to_int501_t(x : std_logic_vector) return int501_t;
subtype uint502_t is unsigned(501 downto 0);
constant uint502_t_SLV_LEN : integer := 502;
function uint502_t_to_slv(x : uint502_t) return std_logic_vector;
function slv_to_uint502_t(x : std_logic_vector) return uint502_t;
subtype int502_t is signed(501 downto 0);
constant int502_t_SLV_LEN : integer := 502;
function int502_t_to_slv(x : int502_t) return std_logic_vector;
function slv_to_int502_t(x : std_logic_vector) return int502_t;
subtype uint503_t is unsigned(502 downto 0);
constant uint503_t_SLV_LEN : integer := 503;
function uint503_t_to_slv(x : uint503_t) return std_logic_vector;
function slv_to_uint503_t(x : std_logic_vector) return uint503_t;
subtype int503_t is signed(502 downto 0);
constant int503_t_SLV_LEN : integer := 503;
function int503_t_to_slv(x : int503_t) return std_logic_vector;
function slv_to_int503_t(x : std_logic_vector) return int503_t;
subtype uint504_t is unsigned(503 downto 0);
constant uint504_t_SLV_LEN : integer := 504;
function uint504_t_to_slv(x : uint504_t) return std_logic_vector;
function slv_to_uint504_t(x : std_logic_vector) return uint504_t;
subtype int504_t is signed(503 downto 0);
constant int504_t_SLV_LEN : integer := 504;
function int504_t_to_slv(x : int504_t) return std_logic_vector;
function slv_to_int504_t(x : std_logic_vector) return int504_t;
subtype uint505_t is unsigned(504 downto 0);
constant uint505_t_SLV_LEN : integer := 505;
function uint505_t_to_slv(x : uint505_t) return std_logic_vector;
function slv_to_uint505_t(x : std_logic_vector) return uint505_t;
subtype int505_t is signed(504 downto 0);
constant int505_t_SLV_LEN : integer := 505;
function int505_t_to_slv(x : int505_t) return std_logic_vector;
function slv_to_int505_t(x : std_logic_vector) return int505_t;
subtype uint506_t is unsigned(505 downto 0);
constant uint506_t_SLV_LEN : integer := 506;
function uint506_t_to_slv(x : uint506_t) return std_logic_vector;
function slv_to_uint506_t(x : std_logic_vector) return uint506_t;
subtype int506_t is signed(505 downto 0);
constant int506_t_SLV_LEN : integer := 506;
function int506_t_to_slv(x : int506_t) return std_logic_vector;
function slv_to_int506_t(x : std_logic_vector) return int506_t;
subtype uint507_t is unsigned(506 downto 0);
constant uint507_t_SLV_LEN : integer := 507;
function uint507_t_to_slv(x : uint507_t) return std_logic_vector;
function slv_to_uint507_t(x : std_logic_vector) return uint507_t;
subtype int507_t is signed(506 downto 0);
constant int507_t_SLV_LEN : integer := 507;
function int507_t_to_slv(x : int507_t) return std_logic_vector;
function slv_to_int507_t(x : std_logic_vector) return int507_t;
subtype uint508_t is unsigned(507 downto 0);
constant uint508_t_SLV_LEN : integer := 508;
function uint508_t_to_slv(x : uint508_t) return std_logic_vector;
function slv_to_uint508_t(x : std_logic_vector) return uint508_t;
subtype int508_t is signed(507 downto 0);
constant int508_t_SLV_LEN : integer := 508;
function int508_t_to_slv(x : int508_t) return std_logic_vector;
function slv_to_int508_t(x : std_logic_vector) return int508_t;
subtype uint509_t is unsigned(508 downto 0);
constant uint509_t_SLV_LEN : integer := 509;
function uint509_t_to_slv(x : uint509_t) return std_logic_vector;
function slv_to_uint509_t(x : std_logic_vector) return uint509_t;
subtype int509_t is signed(508 downto 0);
constant int509_t_SLV_LEN : integer := 509;
function int509_t_to_slv(x : int509_t) return std_logic_vector;
function slv_to_int509_t(x : std_logic_vector) return int509_t;
subtype uint510_t is unsigned(509 downto 0);
constant uint510_t_SLV_LEN : integer := 510;
function uint510_t_to_slv(x : uint510_t) return std_logic_vector;
function slv_to_uint510_t(x : std_logic_vector) return uint510_t;
subtype int510_t is signed(509 downto 0);
constant int510_t_SLV_LEN : integer := 510;
function int510_t_to_slv(x : int510_t) return std_logic_vector;
function slv_to_int510_t(x : std_logic_vector) return int510_t;
subtype uint511_t is unsigned(510 downto 0);
constant uint511_t_SLV_LEN : integer := 511;
function uint511_t_to_slv(x : uint511_t) return std_logic_vector;
function slv_to_uint511_t(x : std_logic_vector) return uint511_t;
subtype int511_t is signed(510 downto 0);
constant int511_t_SLV_LEN : integer := 511;
function int511_t_to_slv(x : int511_t) return std_logic_vector;
function slv_to_int511_t(x : std_logic_vector) return int511_t;
subtype uint512_t is unsigned(511 downto 0);
constant uint512_t_SLV_LEN : integer := 512;
function uint512_t_to_slv(x : uint512_t) return std_logic_vector;
function slv_to_uint512_t(x : std_logic_vector) return uint512_t;
subtype int512_t is signed(511 downto 0);
constant int512_t_SLV_LEN : integer := 512;
function int512_t_to_slv(x : int512_t) return std_logic_vector;
function slv_to_int512_t(x : std_logic_vector) return int512_t;
subtype uint513_t is unsigned(512 downto 0);
constant uint513_t_SLV_LEN : integer := 513;
function uint513_t_to_slv(x : uint513_t) return std_logic_vector;
function slv_to_uint513_t(x : std_logic_vector) return uint513_t;
subtype int513_t is signed(512 downto 0);
constant int513_t_SLV_LEN : integer := 513;
function int513_t_to_slv(x : int513_t) return std_logic_vector;
function slv_to_int513_t(x : std_logic_vector) return int513_t;
subtype uint514_t is unsigned(513 downto 0);
constant uint514_t_SLV_LEN : integer := 514;
function uint514_t_to_slv(x : uint514_t) return std_logic_vector;
function slv_to_uint514_t(x : std_logic_vector) return uint514_t;
subtype int514_t is signed(513 downto 0);
constant int514_t_SLV_LEN : integer := 514;
function int514_t_to_slv(x : int514_t) return std_logic_vector;
function slv_to_int514_t(x : std_logic_vector) return int514_t;
subtype uint515_t is unsigned(514 downto 0);
constant uint515_t_SLV_LEN : integer := 515;
function uint515_t_to_slv(x : uint515_t) return std_logic_vector;
function slv_to_uint515_t(x : std_logic_vector) return uint515_t;
subtype int515_t is signed(514 downto 0);
constant int515_t_SLV_LEN : integer := 515;
function int515_t_to_slv(x : int515_t) return std_logic_vector;
function slv_to_int515_t(x : std_logic_vector) return int515_t;
subtype uint516_t is unsigned(515 downto 0);
constant uint516_t_SLV_LEN : integer := 516;
function uint516_t_to_slv(x : uint516_t) return std_logic_vector;
function slv_to_uint516_t(x : std_logic_vector) return uint516_t;
subtype int516_t is signed(515 downto 0);
constant int516_t_SLV_LEN : integer := 516;
function int516_t_to_slv(x : int516_t) return std_logic_vector;
function slv_to_int516_t(x : std_logic_vector) return int516_t;
subtype uint517_t is unsigned(516 downto 0);
constant uint517_t_SLV_LEN : integer := 517;
function uint517_t_to_slv(x : uint517_t) return std_logic_vector;
function slv_to_uint517_t(x : std_logic_vector) return uint517_t;
subtype int517_t is signed(516 downto 0);
constant int517_t_SLV_LEN : integer := 517;
function int517_t_to_slv(x : int517_t) return std_logic_vector;
function slv_to_int517_t(x : std_logic_vector) return int517_t;
subtype uint518_t is unsigned(517 downto 0);
constant uint518_t_SLV_LEN : integer := 518;
function uint518_t_to_slv(x : uint518_t) return std_logic_vector;
function slv_to_uint518_t(x : std_logic_vector) return uint518_t;
subtype int518_t is signed(517 downto 0);
constant int518_t_SLV_LEN : integer := 518;
function int518_t_to_slv(x : int518_t) return std_logic_vector;
function slv_to_int518_t(x : std_logic_vector) return int518_t;
subtype uint519_t is unsigned(518 downto 0);
constant uint519_t_SLV_LEN : integer := 519;
function uint519_t_to_slv(x : uint519_t) return std_logic_vector;
function slv_to_uint519_t(x : std_logic_vector) return uint519_t;
subtype int519_t is signed(518 downto 0);
constant int519_t_SLV_LEN : integer := 519;
function int519_t_to_slv(x : int519_t) return std_logic_vector;
function slv_to_int519_t(x : std_logic_vector) return int519_t;
subtype uint520_t is unsigned(519 downto 0);
constant uint520_t_SLV_LEN : integer := 520;
function uint520_t_to_slv(x : uint520_t) return std_logic_vector;
function slv_to_uint520_t(x : std_logic_vector) return uint520_t;
subtype int520_t is signed(519 downto 0);
constant int520_t_SLV_LEN : integer := 520;
function int520_t_to_slv(x : int520_t) return std_logic_vector;
function slv_to_int520_t(x : std_logic_vector) return int520_t;
subtype uint521_t is unsigned(520 downto 0);
constant uint521_t_SLV_LEN : integer := 521;
function uint521_t_to_slv(x : uint521_t) return std_logic_vector;
function slv_to_uint521_t(x : std_logic_vector) return uint521_t;
subtype int521_t is signed(520 downto 0);
constant int521_t_SLV_LEN : integer := 521;
function int521_t_to_slv(x : int521_t) return std_logic_vector;
function slv_to_int521_t(x : std_logic_vector) return int521_t;
subtype uint522_t is unsigned(521 downto 0);
constant uint522_t_SLV_LEN : integer := 522;
function uint522_t_to_slv(x : uint522_t) return std_logic_vector;
function slv_to_uint522_t(x : std_logic_vector) return uint522_t;
subtype int522_t is signed(521 downto 0);
constant int522_t_SLV_LEN : integer := 522;
function int522_t_to_slv(x : int522_t) return std_logic_vector;
function slv_to_int522_t(x : std_logic_vector) return int522_t;
subtype uint523_t is unsigned(522 downto 0);
constant uint523_t_SLV_LEN : integer := 523;
function uint523_t_to_slv(x : uint523_t) return std_logic_vector;
function slv_to_uint523_t(x : std_logic_vector) return uint523_t;
subtype int523_t is signed(522 downto 0);
constant int523_t_SLV_LEN : integer := 523;
function int523_t_to_slv(x : int523_t) return std_logic_vector;
function slv_to_int523_t(x : std_logic_vector) return int523_t;
subtype uint524_t is unsigned(523 downto 0);
constant uint524_t_SLV_LEN : integer := 524;
function uint524_t_to_slv(x : uint524_t) return std_logic_vector;
function slv_to_uint524_t(x : std_logic_vector) return uint524_t;
subtype int524_t is signed(523 downto 0);
constant int524_t_SLV_LEN : integer := 524;
function int524_t_to_slv(x : int524_t) return std_logic_vector;
function slv_to_int524_t(x : std_logic_vector) return int524_t;
subtype uint525_t is unsigned(524 downto 0);
constant uint525_t_SLV_LEN : integer := 525;
function uint525_t_to_slv(x : uint525_t) return std_logic_vector;
function slv_to_uint525_t(x : std_logic_vector) return uint525_t;
subtype int525_t is signed(524 downto 0);
constant int525_t_SLV_LEN : integer := 525;
function int525_t_to_slv(x : int525_t) return std_logic_vector;
function slv_to_int525_t(x : std_logic_vector) return int525_t;
subtype uint526_t is unsigned(525 downto 0);
constant uint526_t_SLV_LEN : integer := 526;
function uint526_t_to_slv(x : uint526_t) return std_logic_vector;
function slv_to_uint526_t(x : std_logic_vector) return uint526_t;
subtype int526_t is signed(525 downto 0);
constant int526_t_SLV_LEN : integer := 526;
function int526_t_to_slv(x : int526_t) return std_logic_vector;
function slv_to_int526_t(x : std_logic_vector) return int526_t;
subtype uint527_t is unsigned(526 downto 0);
constant uint527_t_SLV_LEN : integer := 527;
function uint527_t_to_slv(x : uint527_t) return std_logic_vector;
function slv_to_uint527_t(x : std_logic_vector) return uint527_t;
subtype int527_t is signed(526 downto 0);
constant int527_t_SLV_LEN : integer := 527;
function int527_t_to_slv(x : int527_t) return std_logic_vector;
function slv_to_int527_t(x : std_logic_vector) return int527_t;
subtype uint528_t is unsigned(527 downto 0);
constant uint528_t_SLV_LEN : integer := 528;
function uint528_t_to_slv(x : uint528_t) return std_logic_vector;
function slv_to_uint528_t(x : std_logic_vector) return uint528_t;
subtype int528_t is signed(527 downto 0);
constant int528_t_SLV_LEN : integer := 528;
function int528_t_to_slv(x : int528_t) return std_logic_vector;
function slv_to_int528_t(x : std_logic_vector) return int528_t;
subtype uint529_t is unsigned(528 downto 0);
constant uint529_t_SLV_LEN : integer := 529;
function uint529_t_to_slv(x : uint529_t) return std_logic_vector;
function slv_to_uint529_t(x : std_logic_vector) return uint529_t;
subtype int529_t is signed(528 downto 0);
constant int529_t_SLV_LEN : integer := 529;
function int529_t_to_slv(x : int529_t) return std_logic_vector;
function slv_to_int529_t(x : std_logic_vector) return int529_t;
subtype uint530_t is unsigned(529 downto 0);
constant uint530_t_SLV_LEN : integer := 530;
function uint530_t_to_slv(x : uint530_t) return std_logic_vector;
function slv_to_uint530_t(x : std_logic_vector) return uint530_t;
subtype int530_t is signed(529 downto 0);
constant int530_t_SLV_LEN : integer := 530;
function int530_t_to_slv(x : int530_t) return std_logic_vector;
function slv_to_int530_t(x : std_logic_vector) return int530_t;
subtype uint531_t is unsigned(530 downto 0);
constant uint531_t_SLV_LEN : integer := 531;
function uint531_t_to_slv(x : uint531_t) return std_logic_vector;
function slv_to_uint531_t(x : std_logic_vector) return uint531_t;
subtype int531_t is signed(530 downto 0);
constant int531_t_SLV_LEN : integer := 531;
function int531_t_to_slv(x : int531_t) return std_logic_vector;
function slv_to_int531_t(x : std_logic_vector) return int531_t;
subtype uint532_t is unsigned(531 downto 0);
constant uint532_t_SLV_LEN : integer := 532;
function uint532_t_to_slv(x : uint532_t) return std_logic_vector;
function slv_to_uint532_t(x : std_logic_vector) return uint532_t;
subtype int532_t is signed(531 downto 0);
constant int532_t_SLV_LEN : integer := 532;
function int532_t_to_slv(x : int532_t) return std_logic_vector;
function slv_to_int532_t(x : std_logic_vector) return int532_t;
subtype uint533_t is unsigned(532 downto 0);
constant uint533_t_SLV_LEN : integer := 533;
function uint533_t_to_slv(x : uint533_t) return std_logic_vector;
function slv_to_uint533_t(x : std_logic_vector) return uint533_t;
subtype int533_t is signed(532 downto 0);
constant int533_t_SLV_LEN : integer := 533;
function int533_t_to_slv(x : int533_t) return std_logic_vector;
function slv_to_int533_t(x : std_logic_vector) return int533_t;
subtype uint534_t is unsigned(533 downto 0);
constant uint534_t_SLV_LEN : integer := 534;
function uint534_t_to_slv(x : uint534_t) return std_logic_vector;
function slv_to_uint534_t(x : std_logic_vector) return uint534_t;
subtype int534_t is signed(533 downto 0);
constant int534_t_SLV_LEN : integer := 534;
function int534_t_to_slv(x : int534_t) return std_logic_vector;
function slv_to_int534_t(x : std_logic_vector) return int534_t;
subtype uint535_t is unsigned(534 downto 0);
constant uint535_t_SLV_LEN : integer := 535;
function uint535_t_to_slv(x : uint535_t) return std_logic_vector;
function slv_to_uint535_t(x : std_logic_vector) return uint535_t;
subtype int535_t is signed(534 downto 0);
constant int535_t_SLV_LEN : integer := 535;
function int535_t_to_slv(x : int535_t) return std_logic_vector;
function slv_to_int535_t(x : std_logic_vector) return int535_t;
subtype uint536_t is unsigned(535 downto 0);
constant uint536_t_SLV_LEN : integer := 536;
function uint536_t_to_slv(x : uint536_t) return std_logic_vector;
function slv_to_uint536_t(x : std_logic_vector) return uint536_t;
subtype int536_t is signed(535 downto 0);
constant int536_t_SLV_LEN : integer := 536;
function int536_t_to_slv(x : int536_t) return std_logic_vector;
function slv_to_int536_t(x : std_logic_vector) return int536_t;
subtype uint537_t is unsigned(536 downto 0);
constant uint537_t_SLV_LEN : integer := 537;
function uint537_t_to_slv(x : uint537_t) return std_logic_vector;
function slv_to_uint537_t(x : std_logic_vector) return uint537_t;
subtype int537_t is signed(536 downto 0);
constant int537_t_SLV_LEN : integer := 537;
function int537_t_to_slv(x : int537_t) return std_logic_vector;
function slv_to_int537_t(x : std_logic_vector) return int537_t;
subtype uint538_t is unsigned(537 downto 0);
constant uint538_t_SLV_LEN : integer := 538;
function uint538_t_to_slv(x : uint538_t) return std_logic_vector;
function slv_to_uint538_t(x : std_logic_vector) return uint538_t;
subtype int538_t is signed(537 downto 0);
constant int538_t_SLV_LEN : integer := 538;
function int538_t_to_slv(x : int538_t) return std_logic_vector;
function slv_to_int538_t(x : std_logic_vector) return int538_t;
subtype uint539_t is unsigned(538 downto 0);
constant uint539_t_SLV_LEN : integer := 539;
function uint539_t_to_slv(x : uint539_t) return std_logic_vector;
function slv_to_uint539_t(x : std_logic_vector) return uint539_t;
subtype int539_t is signed(538 downto 0);
constant int539_t_SLV_LEN : integer := 539;
function int539_t_to_slv(x : int539_t) return std_logic_vector;
function slv_to_int539_t(x : std_logic_vector) return int539_t;
subtype uint540_t is unsigned(539 downto 0);
constant uint540_t_SLV_LEN : integer := 540;
function uint540_t_to_slv(x : uint540_t) return std_logic_vector;
function slv_to_uint540_t(x : std_logic_vector) return uint540_t;
subtype int540_t is signed(539 downto 0);
constant int540_t_SLV_LEN : integer := 540;
function int540_t_to_slv(x : int540_t) return std_logic_vector;
function slv_to_int540_t(x : std_logic_vector) return int540_t;
subtype uint541_t is unsigned(540 downto 0);
constant uint541_t_SLV_LEN : integer := 541;
function uint541_t_to_slv(x : uint541_t) return std_logic_vector;
function slv_to_uint541_t(x : std_logic_vector) return uint541_t;
subtype int541_t is signed(540 downto 0);
constant int541_t_SLV_LEN : integer := 541;
function int541_t_to_slv(x : int541_t) return std_logic_vector;
function slv_to_int541_t(x : std_logic_vector) return int541_t;
subtype uint542_t is unsigned(541 downto 0);
constant uint542_t_SLV_LEN : integer := 542;
function uint542_t_to_slv(x : uint542_t) return std_logic_vector;
function slv_to_uint542_t(x : std_logic_vector) return uint542_t;
subtype int542_t is signed(541 downto 0);
constant int542_t_SLV_LEN : integer := 542;
function int542_t_to_slv(x : int542_t) return std_logic_vector;
function slv_to_int542_t(x : std_logic_vector) return int542_t;
subtype uint543_t is unsigned(542 downto 0);
constant uint543_t_SLV_LEN : integer := 543;
function uint543_t_to_slv(x : uint543_t) return std_logic_vector;
function slv_to_uint543_t(x : std_logic_vector) return uint543_t;
subtype int543_t is signed(542 downto 0);
constant int543_t_SLV_LEN : integer := 543;
function int543_t_to_slv(x : int543_t) return std_logic_vector;
function slv_to_int543_t(x : std_logic_vector) return int543_t;
subtype uint544_t is unsigned(543 downto 0);
constant uint544_t_SLV_LEN : integer := 544;
function uint544_t_to_slv(x : uint544_t) return std_logic_vector;
function slv_to_uint544_t(x : std_logic_vector) return uint544_t;
subtype int544_t is signed(543 downto 0);
constant int544_t_SLV_LEN : integer := 544;
function int544_t_to_slv(x : int544_t) return std_logic_vector;
function slv_to_int544_t(x : std_logic_vector) return int544_t;
subtype uint545_t is unsigned(544 downto 0);
constant uint545_t_SLV_LEN : integer := 545;
function uint545_t_to_slv(x : uint545_t) return std_logic_vector;
function slv_to_uint545_t(x : std_logic_vector) return uint545_t;
subtype int545_t is signed(544 downto 0);
constant int545_t_SLV_LEN : integer := 545;
function int545_t_to_slv(x : int545_t) return std_logic_vector;
function slv_to_int545_t(x : std_logic_vector) return int545_t;
subtype uint546_t is unsigned(545 downto 0);
constant uint546_t_SLV_LEN : integer := 546;
function uint546_t_to_slv(x : uint546_t) return std_logic_vector;
function slv_to_uint546_t(x : std_logic_vector) return uint546_t;
subtype int546_t is signed(545 downto 0);
constant int546_t_SLV_LEN : integer := 546;
function int546_t_to_slv(x : int546_t) return std_logic_vector;
function slv_to_int546_t(x : std_logic_vector) return int546_t;
subtype uint547_t is unsigned(546 downto 0);
constant uint547_t_SLV_LEN : integer := 547;
function uint547_t_to_slv(x : uint547_t) return std_logic_vector;
function slv_to_uint547_t(x : std_logic_vector) return uint547_t;
subtype int547_t is signed(546 downto 0);
constant int547_t_SLV_LEN : integer := 547;
function int547_t_to_slv(x : int547_t) return std_logic_vector;
function slv_to_int547_t(x : std_logic_vector) return int547_t;
subtype uint548_t is unsigned(547 downto 0);
constant uint548_t_SLV_LEN : integer := 548;
function uint548_t_to_slv(x : uint548_t) return std_logic_vector;
function slv_to_uint548_t(x : std_logic_vector) return uint548_t;
subtype int548_t is signed(547 downto 0);
constant int548_t_SLV_LEN : integer := 548;
function int548_t_to_slv(x : int548_t) return std_logic_vector;
function slv_to_int548_t(x : std_logic_vector) return int548_t;
subtype uint549_t is unsigned(548 downto 0);
constant uint549_t_SLV_LEN : integer := 549;
function uint549_t_to_slv(x : uint549_t) return std_logic_vector;
function slv_to_uint549_t(x : std_logic_vector) return uint549_t;
subtype int549_t is signed(548 downto 0);
constant int549_t_SLV_LEN : integer := 549;
function int549_t_to_slv(x : int549_t) return std_logic_vector;
function slv_to_int549_t(x : std_logic_vector) return int549_t;
subtype uint550_t is unsigned(549 downto 0);
constant uint550_t_SLV_LEN : integer := 550;
function uint550_t_to_slv(x : uint550_t) return std_logic_vector;
function slv_to_uint550_t(x : std_logic_vector) return uint550_t;
subtype int550_t is signed(549 downto 0);
constant int550_t_SLV_LEN : integer := 550;
function int550_t_to_slv(x : int550_t) return std_logic_vector;
function slv_to_int550_t(x : std_logic_vector) return int550_t;
subtype uint551_t is unsigned(550 downto 0);
constant uint551_t_SLV_LEN : integer := 551;
function uint551_t_to_slv(x : uint551_t) return std_logic_vector;
function slv_to_uint551_t(x : std_logic_vector) return uint551_t;
subtype int551_t is signed(550 downto 0);
constant int551_t_SLV_LEN : integer := 551;
function int551_t_to_slv(x : int551_t) return std_logic_vector;
function slv_to_int551_t(x : std_logic_vector) return int551_t;
subtype uint552_t is unsigned(551 downto 0);
constant uint552_t_SLV_LEN : integer := 552;
function uint552_t_to_slv(x : uint552_t) return std_logic_vector;
function slv_to_uint552_t(x : std_logic_vector) return uint552_t;
subtype int552_t is signed(551 downto 0);
constant int552_t_SLV_LEN : integer := 552;
function int552_t_to_slv(x : int552_t) return std_logic_vector;
function slv_to_int552_t(x : std_logic_vector) return int552_t;
subtype uint553_t is unsigned(552 downto 0);
constant uint553_t_SLV_LEN : integer := 553;
function uint553_t_to_slv(x : uint553_t) return std_logic_vector;
function slv_to_uint553_t(x : std_logic_vector) return uint553_t;
subtype int553_t is signed(552 downto 0);
constant int553_t_SLV_LEN : integer := 553;
function int553_t_to_slv(x : int553_t) return std_logic_vector;
function slv_to_int553_t(x : std_logic_vector) return int553_t;
subtype uint554_t is unsigned(553 downto 0);
constant uint554_t_SLV_LEN : integer := 554;
function uint554_t_to_slv(x : uint554_t) return std_logic_vector;
function slv_to_uint554_t(x : std_logic_vector) return uint554_t;
subtype int554_t is signed(553 downto 0);
constant int554_t_SLV_LEN : integer := 554;
function int554_t_to_slv(x : int554_t) return std_logic_vector;
function slv_to_int554_t(x : std_logic_vector) return int554_t;
subtype uint555_t is unsigned(554 downto 0);
constant uint555_t_SLV_LEN : integer := 555;
function uint555_t_to_slv(x : uint555_t) return std_logic_vector;
function slv_to_uint555_t(x : std_logic_vector) return uint555_t;
subtype int555_t is signed(554 downto 0);
constant int555_t_SLV_LEN : integer := 555;
function int555_t_to_slv(x : int555_t) return std_logic_vector;
function slv_to_int555_t(x : std_logic_vector) return int555_t;
subtype uint556_t is unsigned(555 downto 0);
constant uint556_t_SLV_LEN : integer := 556;
function uint556_t_to_slv(x : uint556_t) return std_logic_vector;
function slv_to_uint556_t(x : std_logic_vector) return uint556_t;
subtype int556_t is signed(555 downto 0);
constant int556_t_SLV_LEN : integer := 556;
function int556_t_to_slv(x : int556_t) return std_logic_vector;
function slv_to_int556_t(x : std_logic_vector) return int556_t;
subtype uint557_t is unsigned(556 downto 0);
constant uint557_t_SLV_LEN : integer := 557;
function uint557_t_to_slv(x : uint557_t) return std_logic_vector;
function slv_to_uint557_t(x : std_logic_vector) return uint557_t;
subtype int557_t is signed(556 downto 0);
constant int557_t_SLV_LEN : integer := 557;
function int557_t_to_slv(x : int557_t) return std_logic_vector;
function slv_to_int557_t(x : std_logic_vector) return int557_t;
subtype uint558_t is unsigned(557 downto 0);
constant uint558_t_SLV_LEN : integer := 558;
function uint558_t_to_slv(x : uint558_t) return std_logic_vector;
function slv_to_uint558_t(x : std_logic_vector) return uint558_t;
subtype int558_t is signed(557 downto 0);
constant int558_t_SLV_LEN : integer := 558;
function int558_t_to_slv(x : int558_t) return std_logic_vector;
function slv_to_int558_t(x : std_logic_vector) return int558_t;
subtype uint559_t is unsigned(558 downto 0);
constant uint559_t_SLV_LEN : integer := 559;
function uint559_t_to_slv(x : uint559_t) return std_logic_vector;
function slv_to_uint559_t(x : std_logic_vector) return uint559_t;
subtype int559_t is signed(558 downto 0);
constant int559_t_SLV_LEN : integer := 559;
function int559_t_to_slv(x : int559_t) return std_logic_vector;
function slv_to_int559_t(x : std_logic_vector) return int559_t;
subtype uint560_t is unsigned(559 downto 0);
constant uint560_t_SLV_LEN : integer := 560;
function uint560_t_to_slv(x : uint560_t) return std_logic_vector;
function slv_to_uint560_t(x : std_logic_vector) return uint560_t;
subtype int560_t is signed(559 downto 0);
constant int560_t_SLV_LEN : integer := 560;
function int560_t_to_slv(x : int560_t) return std_logic_vector;
function slv_to_int560_t(x : std_logic_vector) return int560_t;
subtype uint561_t is unsigned(560 downto 0);
constant uint561_t_SLV_LEN : integer := 561;
function uint561_t_to_slv(x : uint561_t) return std_logic_vector;
function slv_to_uint561_t(x : std_logic_vector) return uint561_t;
subtype int561_t is signed(560 downto 0);
constant int561_t_SLV_LEN : integer := 561;
function int561_t_to_slv(x : int561_t) return std_logic_vector;
function slv_to_int561_t(x : std_logic_vector) return int561_t;
subtype uint562_t is unsigned(561 downto 0);
constant uint562_t_SLV_LEN : integer := 562;
function uint562_t_to_slv(x : uint562_t) return std_logic_vector;
function slv_to_uint562_t(x : std_logic_vector) return uint562_t;
subtype int562_t is signed(561 downto 0);
constant int562_t_SLV_LEN : integer := 562;
function int562_t_to_slv(x : int562_t) return std_logic_vector;
function slv_to_int562_t(x : std_logic_vector) return int562_t;
subtype uint563_t is unsigned(562 downto 0);
constant uint563_t_SLV_LEN : integer := 563;
function uint563_t_to_slv(x : uint563_t) return std_logic_vector;
function slv_to_uint563_t(x : std_logic_vector) return uint563_t;
subtype int563_t is signed(562 downto 0);
constant int563_t_SLV_LEN : integer := 563;
function int563_t_to_slv(x : int563_t) return std_logic_vector;
function slv_to_int563_t(x : std_logic_vector) return int563_t;
subtype uint564_t is unsigned(563 downto 0);
constant uint564_t_SLV_LEN : integer := 564;
function uint564_t_to_slv(x : uint564_t) return std_logic_vector;
function slv_to_uint564_t(x : std_logic_vector) return uint564_t;
subtype int564_t is signed(563 downto 0);
constant int564_t_SLV_LEN : integer := 564;
function int564_t_to_slv(x : int564_t) return std_logic_vector;
function slv_to_int564_t(x : std_logic_vector) return int564_t;
subtype uint565_t is unsigned(564 downto 0);
constant uint565_t_SLV_LEN : integer := 565;
function uint565_t_to_slv(x : uint565_t) return std_logic_vector;
function slv_to_uint565_t(x : std_logic_vector) return uint565_t;
subtype int565_t is signed(564 downto 0);
constant int565_t_SLV_LEN : integer := 565;
function int565_t_to_slv(x : int565_t) return std_logic_vector;
function slv_to_int565_t(x : std_logic_vector) return int565_t;
subtype uint566_t is unsigned(565 downto 0);
constant uint566_t_SLV_LEN : integer := 566;
function uint566_t_to_slv(x : uint566_t) return std_logic_vector;
function slv_to_uint566_t(x : std_logic_vector) return uint566_t;
subtype int566_t is signed(565 downto 0);
constant int566_t_SLV_LEN : integer := 566;
function int566_t_to_slv(x : int566_t) return std_logic_vector;
function slv_to_int566_t(x : std_logic_vector) return int566_t;
subtype uint567_t is unsigned(566 downto 0);
constant uint567_t_SLV_LEN : integer := 567;
function uint567_t_to_slv(x : uint567_t) return std_logic_vector;
function slv_to_uint567_t(x : std_logic_vector) return uint567_t;
subtype int567_t is signed(566 downto 0);
constant int567_t_SLV_LEN : integer := 567;
function int567_t_to_slv(x : int567_t) return std_logic_vector;
function slv_to_int567_t(x : std_logic_vector) return int567_t;
subtype uint568_t is unsigned(567 downto 0);
constant uint568_t_SLV_LEN : integer := 568;
function uint568_t_to_slv(x : uint568_t) return std_logic_vector;
function slv_to_uint568_t(x : std_logic_vector) return uint568_t;
subtype int568_t is signed(567 downto 0);
constant int568_t_SLV_LEN : integer := 568;
function int568_t_to_slv(x : int568_t) return std_logic_vector;
function slv_to_int568_t(x : std_logic_vector) return int568_t;
subtype uint569_t is unsigned(568 downto 0);
constant uint569_t_SLV_LEN : integer := 569;
function uint569_t_to_slv(x : uint569_t) return std_logic_vector;
function slv_to_uint569_t(x : std_logic_vector) return uint569_t;
subtype int569_t is signed(568 downto 0);
constant int569_t_SLV_LEN : integer := 569;
function int569_t_to_slv(x : int569_t) return std_logic_vector;
function slv_to_int569_t(x : std_logic_vector) return int569_t;
subtype uint570_t is unsigned(569 downto 0);
constant uint570_t_SLV_LEN : integer := 570;
function uint570_t_to_slv(x : uint570_t) return std_logic_vector;
function slv_to_uint570_t(x : std_logic_vector) return uint570_t;
subtype int570_t is signed(569 downto 0);
constant int570_t_SLV_LEN : integer := 570;
function int570_t_to_slv(x : int570_t) return std_logic_vector;
function slv_to_int570_t(x : std_logic_vector) return int570_t;
subtype uint571_t is unsigned(570 downto 0);
constant uint571_t_SLV_LEN : integer := 571;
function uint571_t_to_slv(x : uint571_t) return std_logic_vector;
function slv_to_uint571_t(x : std_logic_vector) return uint571_t;
subtype int571_t is signed(570 downto 0);
constant int571_t_SLV_LEN : integer := 571;
function int571_t_to_slv(x : int571_t) return std_logic_vector;
function slv_to_int571_t(x : std_logic_vector) return int571_t;
subtype uint572_t is unsigned(571 downto 0);
constant uint572_t_SLV_LEN : integer := 572;
function uint572_t_to_slv(x : uint572_t) return std_logic_vector;
function slv_to_uint572_t(x : std_logic_vector) return uint572_t;
subtype int572_t is signed(571 downto 0);
constant int572_t_SLV_LEN : integer := 572;
function int572_t_to_slv(x : int572_t) return std_logic_vector;
function slv_to_int572_t(x : std_logic_vector) return int572_t;
subtype uint573_t is unsigned(572 downto 0);
constant uint573_t_SLV_LEN : integer := 573;
function uint573_t_to_slv(x : uint573_t) return std_logic_vector;
function slv_to_uint573_t(x : std_logic_vector) return uint573_t;
subtype int573_t is signed(572 downto 0);
constant int573_t_SLV_LEN : integer := 573;
function int573_t_to_slv(x : int573_t) return std_logic_vector;
function slv_to_int573_t(x : std_logic_vector) return int573_t;
subtype uint574_t is unsigned(573 downto 0);
constant uint574_t_SLV_LEN : integer := 574;
function uint574_t_to_slv(x : uint574_t) return std_logic_vector;
function slv_to_uint574_t(x : std_logic_vector) return uint574_t;
subtype int574_t is signed(573 downto 0);
constant int574_t_SLV_LEN : integer := 574;
function int574_t_to_slv(x : int574_t) return std_logic_vector;
function slv_to_int574_t(x : std_logic_vector) return int574_t;
subtype uint575_t is unsigned(574 downto 0);
constant uint575_t_SLV_LEN : integer := 575;
function uint575_t_to_slv(x : uint575_t) return std_logic_vector;
function slv_to_uint575_t(x : std_logic_vector) return uint575_t;
subtype int575_t is signed(574 downto 0);
constant int575_t_SLV_LEN : integer := 575;
function int575_t_to_slv(x : int575_t) return std_logic_vector;
function slv_to_int575_t(x : std_logic_vector) return int575_t;
subtype uint576_t is unsigned(575 downto 0);
constant uint576_t_SLV_LEN : integer := 576;
function uint576_t_to_slv(x : uint576_t) return std_logic_vector;
function slv_to_uint576_t(x : std_logic_vector) return uint576_t;
subtype int576_t is signed(575 downto 0);
constant int576_t_SLV_LEN : integer := 576;
function int576_t_to_slv(x : int576_t) return std_logic_vector;
function slv_to_int576_t(x : std_logic_vector) return int576_t;
subtype uint577_t is unsigned(576 downto 0);
constant uint577_t_SLV_LEN : integer := 577;
function uint577_t_to_slv(x : uint577_t) return std_logic_vector;
function slv_to_uint577_t(x : std_logic_vector) return uint577_t;
subtype int577_t is signed(576 downto 0);
constant int577_t_SLV_LEN : integer := 577;
function int577_t_to_slv(x : int577_t) return std_logic_vector;
function slv_to_int577_t(x : std_logic_vector) return int577_t;
subtype uint578_t is unsigned(577 downto 0);
constant uint578_t_SLV_LEN : integer := 578;
function uint578_t_to_slv(x : uint578_t) return std_logic_vector;
function slv_to_uint578_t(x : std_logic_vector) return uint578_t;
subtype int578_t is signed(577 downto 0);
constant int578_t_SLV_LEN : integer := 578;
function int578_t_to_slv(x : int578_t) return std_logic_vector;
function slv_to_int578_t(x : std_logic_vector) return int578_t;
subtype uint579_t is unsigned(578 downto 0);
constant uint579_t_SLV_LEN : integer := 579;
function uint579_t_to_slv(x : uint579_t) return std_logic_vector;
function slv_to_uint579_t(x : std_logic_vector) return uint579_t;
subtype int579_t is signed(578 downto 0);
constant int579_t_SLV_LEN : integer := 579;
function int579_t_to_slv(x : int579_t) return std_logic_vector;
function slv_to_int579_t(x : std_logic_vector) return int579_t;
subtype uint580_t is unsigned(579 downto 0);
constant uint580_t_SLV_LEN : integer := 580;
function uint580_t_to_slv(x : uint580_t) return std_logic_vector;
function slv_to_uint580_t(x : std_logic_vector) return uint580_t;
subtype int580_t is signed(579 downto 0);
constant int580_t_SLV_LEN : integer := 580;
function int580_t_to_slv(x : int580_t) return std_logic_vector;
function slv_to_int580_t(x : std_logic_vector) return int580_t;
subtype uint581_t is unsigned(580 downto 0);
constant uint581_t_SLV_LEN : integer := 581;
function uint581_t_to_slv(x : uint581_t) return std_logic_vector;
function slv_to_uint581_t(x : std_logic_vector) return uint581_t;
subtype int581_t is signed(580 downto 0);
constant int581_t_SLV_LEN : integer := 581;
function int581_t_to_slv(x : int581_t) return std_logic_vector;
function slv_to_int581_t(x : std_logic_vector) return int581_t;
subtype uint582_t is unsigned(581 downto 0);
constant uint582_t_SLV_LEN : integer := 582;
function uint582_t_to_slv(x : uint582_t) return std_logic_vector;
function slv_to_uint582_t(x : std_logic_vector) return uint582_t;
subtype int582_t is signed(581 downto 0);
constant int582_t_SLV_LEN : integer := 582;
function int582_t_to_slv(x : int582_t) return std_logic_vector;
function slv_to_int582_t(x : std_logic_vector) return int582_t;
subtype uint583_t is unsigned(582 downto 0);
constant uint583_t_SLV_LEN : integer := 583;
function uint583_t_to_slv(x : uint583_t) return std_logic_vector;
function slv_to_uint583_t(x : std_logic_vector) return uint583_t;
subtype int583_t is signed(582 downto 0);
constant int583_t_SLV_LEN : integer := 583;
function int583_t_to_slv(x : int583_t) return std_logic_vector;
function slv_to_int583_t(x : std_logic_vector) return int583_t;
subtype uint584_t is unsigned(583 downto 0);
constant uint584_t_SLV_LEN : integer := 584;
function uint584_t_to_slv(x : uint584_t) return std_logic_vector;
function slv_to_uint584_t(x : std_logic_vector) return uint584_t;
subtype int584_t is signed(583 downto 0);
constant int584_t_SLV_LEN : integer := 584;
function int584_t_to_slv(x : int584_t) return std_logic_vector;
function slv_to_int584_t(x : std_logic_vector) return int584_t;
subtype uint585_t is unsigned(584 downto 0);
constant uint585_t_SLV_LEN : integer := 585;
function uint585_t_to_slv(x : uint585_t) return std_logic_vector;
function slv_to_uint585_t(x : std_logic_vector) return uint585_t;
subtype int585_t is signed(584 downto 0);
constant int585_t_SLV_LEN : integer := 585;
function int585_t_to_slv(x : int585_t) return std_logic_vector;
function slv_to_int585_t(x : std_logic_vector) return int585_t;
subtype uint586_t is unsigned(585 downto 0);
constant uint586_t_SLV_LEN : integer := 586;
function uint586_t_to_slv(x : uint586_t) return std_logic_vector;
function slv_to_uint586_t(x : std_logic_vector) return uint586_t;
subtype int586_t is signed(585 downto 0);
constant int586_t_SLV_LEN : integer := 586;
function int586_t_to_slv(x : int586_t) return std_logic_vector;
function slv_to_int586_t(x : std_logic_vector) return int586_t;
subtype uint587_t is unsigned(586 downto 0);
constant uint587_t_SLV_LEN : integer := 587;
function uint587_t_to_slv(x : uint587_t) return std_logic_vector;
function slv_to_uint587_t(x : std_logic_vector) return uint587_t;
subtype int587_t is signed(586 downto 0);
constant int587_t_SLV_LEN : integer := 587;
function int587_t_to_slv(x : int587_t) return std_logic_vector;
function slv_to_int587_t(x : std_logic_vector) return int587_t;
subtype uint588_t is unsigned(587 downto 0);
constant uint588_t_SLV_LEN : integer := 588;
function uint588_t_to_slv(x : uint588_t) return std_logic_vector;
function slv_to_uint588_t(x : std_logic_vector) return uint588_t;
subtype int588_t is signed(587 downto 0);
constant int588_t_SLV_LEN : integer := 588;
function int588_t_to_slv(x : int588_t) return std_logic_vector;
function slv_to_int588_t(x : std_logic_vector) return int588_t;
subtype uint589_t is unsigned(588 downto 0);
constant uint589_t_SLV_LEN : integer := 589;
function uint589_t_to_slv(x : uint589_t) return std_logic_vector;
function slv_to_uint589_t(x : std_logic_vector) return uint589_t;
subtype int589_t is signed(588 downto 0);
constant int589_t_SLV_LEN : integer := 589;
function int589_t_to_slv(x : int589_t) return std_logic_vector;
function slv_to_int589_t(x : std_logic_vector) return int589_t;
subtype uint590_t is unsigned(589 downto 0);
constant uint590_t_SLV_LEN : integer := 590;
function uint590_t_to_slv(x : uint590_t) return std_logic_vector;
function slv_to_uint590_t(x : std_logic_vector) return uint590_t;
subtype int590_t is signed(589 downto 0);
constant int590_t_SLV_LEN : integer := 590;
function int590_t_to_slv(x : int590_t) return std_logic_vector;
function slv_to_int590_t(x : std_logic_vector) return int590_t;
subtype uint591_t is unsigned(590 downto 0);
constant uint591_t_SLV_LEN : integer := 591;
function uint591_t_to_slv(x : uint591_t) return std_logic_vector;
function slv_to_uint591_t(x : std_logic_vector) return uint591_t;
subtype int591_t is signed(590 downto 0);
constant int591_t_SLV_LEN : integer := 591;
function int591_t_to_slv(x : int591_t) return std_logic_vector;
function slv_to_int591_t(x : std_logic_vector) return int591_t;
subtype uint592_t is unsigned(591 downto 0);
constant uint592_t_SLV_LEN : integer := 592;
function uint592_t_to_slv(x : uint592_t) return std_logic_vector;
function slv_to_uint592_t(x : std_logic_vector) return uint592_t;
subtype int592_t is signed(591 downto 0);
constant int592_t_SLV_LEN : integer := 592;
function int592_t_to_slv(x : int592_t) return std_logic_vector;
function slv_to_int592_t(x : std_logic_vector) return int592_t;
subtype uint593_t is unsigned(592 downto 0);
constant uint593_t_SLV_LEN : integer := 593;
function uint593_t_to_slv(x : uint593_t) return std_logic_vector;
function slv_to_uint593_t(x : std_logic_vector) return uint593_t;
subtype int593_t is signed(592 downto 0);
constant int593_t_SLV_LEN : integer := 593;
function int593_t_to_slv(x : int593_t) return std_logic_vector;
function slv_to_int593_t(x : std_logic_vector) return int593_t;
subtype uint594_t is unsigned(593 downto 0);
constant uint594_t_SLV_LEN : integer := 594;
function uint594_t_to_slv(x : uint594_t) return std_logic_vector;
function slv_to_uint594_t(x : std_logic_vector) return uint594_t;
subtype int594_t is signed(593 downto 0);
constant int594_t_SLV_LEN : integer := 594;
function int594_t_to_slv(x : int594_t) return std_logic_vector;
function slv_to_int594_t(x : std_logic_vector) return int594_t;
subtype uint595_t is unsigned(594 downto 0);
constant uint595_t_SLV_LEN : integer := 595;
function uint595_t_to_slv(x : uint595_t) return std_logic_vector;
function slv_to_uint595_t(x : std_logic_vector) return uint595_t;
subtype int595_t is signed(594 downto 0);
constant int595_t_SLV_LEN : integer := 595;
function int595_t_to_slv(x : int595_t) return std_logic_vector;
function slv_to_int595_t(x : std_logic_vector) return int595_t;
subtype uint596_t is unsigned(595 downto 0);
constant uint596_t_SLV_LEN : integer := 596;
function uint596_t_to_slv(x : uint596_t) return std_logic_vector;
function slv_to_uint596_t(x : std_logic_vector) return uint596_t;
subtype int596_t is signed(595 downto 0);
constant int596_t_SLV_LEN : integer := 596;
function int596_t_to_slv(x : int596_t) return std_logic_vector;
function slv_to_int596_t(x : std_logic_vector) return int596_t;
subtype uint597_t is unsigned(596 downto 0);
constant uint597_t_SLV_LEN : integer := 597;
function uint597_t_to_slv(x : uint597_t) return std_logic_vector;
function slv_to_uint597_t(x : std_logic_vector) return uint597_t;
subtype int597_t is signed(596 downto 0);
constant int597_t_SLV_LEN : integer := 597;
function int597_t_to_slv(x : int597_t) return std_logic_vector;
function slv_to_int597_t(x : std_logic_vector) return int597_t;
subtype uint598_t is unsigned(597 downto 0);
constant uint598_t_SLV_LEN : integer := 598;
function uint598_t_to_slv(x : uint598_t) return std_logic_vector;
function slv_to_uint598_t(x : std_logic_vector) return uint598_t;
subtype int598_t is signed(597 downto 0);
constant int598_t_SLV_LEN : integer := 598;
function int598_t_to_slv(x : int598_t) return std_logic_vector;
function slv_to_int598_t(x : std_logic_vector) return int598_t;
subtype uint599_t is unsigned(598 downto 0);
constant uint599_t_SLV_LEN : integer := 599;
function uint599_t_to_slv(x : uint599_t) return std_logic_vector;
function slv_to_uint599_t(x : std_logic_vector) return uint599_t;
subtype int599_t is signed(598 downto 0);
constant int599_t_SLV_LEN : integer := 599;
function int599_t_to_slv(x : int599_t) return std_logic_vector;
function slv_to_int599_t(x : std_logic_vector) return int599_t;
subtype uint600_t is unsigned(599 downto 0);
constant uint600_t_SLV_LEN : integer := 600;
function uint600_t_to_slv(x : uint600_t) return std_logic_vector;
function slv_to_uint600_t(x : std_logic_vector) return uint600_t;
subtype int600_t is signed(599 downto 0);
constant int600_t_SLV_LEN : integer := 600;
function int600_t_to_slv(x : int600_t) return std_logic_vector;
function slv_to_int600_t(x : std_logic_vector) return int600_t;
subtype uint601_t is unsigned(600 downto 0);
constant uint601_t_SLV_LEN : integer := 601;
function uint601_t_to_slv(x : uint601_t) return std_logic_vector;
function slv_to_uint601_t(x : std_logic_vector) return uint601_t;
subtype int601_t is signed(600 downto 0);
constant int601_t_SLV_LEN : integer := 601;
function int601_t_to_slv(x : int601_t) return std_logic_vector;
function slv_to_int601_t(x : std_logic_vector) return int601_t;
subtype uint602_t is unsigned(601 downto 0);
constant uint602_t_SLV_LEN : integer := 602;
function uint602_t_to_slv(x : uint602_t) return std_logic_vector;
function slv_to_uint602_t(x : std_logic_vector) return uint602_t;
subtype int602_t is signed(601 downto 0);
constant int602_t_SLV_LEN : integer := 602;
function int602_t_to_slv(x : int602_t) return std_logic_vector;
function slv_to_int602_t(x : std_logic_vector) return int602_t;
subtype uint603_t is unsigned(602 downto 0);
constant uint603_t_SLV_LEN : integer := 603;
function uint603_t_to_slv(x : uint603_t) return std_logic_vector;
function slv_to_uint603_t(x : std_logic_vector) return uint603_t;
subtype int603_t is signed(602 downto 0);
constant int603_t_SLV_LEN : integer := 603;
function int603_t_to_slv(x : int603_t) return std_logic_vector;
function slv_to_int603_t(x : std_logic_vector) return int603_t;
subtype uint604_t is unsigned(603 downto 0);
constant uint604_t_SLV_LEN : integer := 604;
function uint604_t_to_slv(x : uint604_t) return std_logic_vector;
function slv_to_uint604_t(x : std_logic_vector) return uint604_t;
subtype int604_t is signed(603 downto 0);
constant int604_t_SLV_LEN : integer := 604;
function int604_t_to_slv(x : int604_t) return std_logic_vector;
function slv_to_int604_t(x : std_logic_vector) return int604_t;
subtype uint605_t is unsigned(604 downto 0);
constant uint605_t_SLV_LEN : integer := 605;
function uint605_t_to_slv(x : uint605_t) return std_logic_vector;
function slv_to_uint605_t(x : std_logic_vector) return uint605_t;
subtype int605_t is signed(604 downto 0);
constant int605_t_SLV_LEN : integer := 605;
function int605_t_to_slv(x : int605_t) return std_logic_vector;
function slv_to_int605_t(x : std_logic_vector) return int605_t;
subtype uint606_t is unsigned(605 downto 0);
constant uint606_t_SLV_LEN : integer := 606;
function uint606_t_to_slv(x : uint606_t) return std_logic_vector;
function slv_to_uint606_t(x : std_logic_vector) return uint606_t;
subtype int606_t is signed(605 downto 0);
constant int606_t_SLV_LEN : integer := 606;
function int606_t_to_slv(x : int606_t) return std_logic_vector;
function slv_to_int606_t(x : std_logic_vector) return int606_t;
subtype uint607_t is unsigned(606 downto 0);
constant uint607_t_SLV_LEN : integer := 607;
function uint607_t_to_slv(x : uint607_t) return std_logic_vector;
function slv_to_uint607_t(x : std_logic_vector) return uint607_t;
subtype int607_t is signed(606 downto 0);
constant int607_t_SLV_LEN : integer := 607;
function int607_t_to_slv(x : int607_t) return std_logic_vector;
function slv_to_int607_t(x : std_logic_vector) return int607_t;
subtype uint608_t is unsigned(607 downto 0);
constant uint608_t_SLV_LEN : integer := 608;
function uint608_t_to_slv(x : uint608_t) return std_logic_vector;
function slv_to_uint608_t(x : std_logic_vector) return uint608_t;
subtype int608_t is signed(607 downto 0);
constant int608_t_SLV_LEN : integer := 608;
function int608_t_to_slv(x : int608_t) return std_logic_vector;
function slv_to_int608_t(x : std_logic_vector) return int608_t;
subtype uint609_t is unsigned(608 downto 0);
constant uint609_t_SLV_LEN : integer := 609;
function uint609_t_to_slv(x : uint609_t) return std_logic_vector;
function slv_to_uint609_t(x : std_logic_vector) return uint609_t;
subtype int609_t is signed(608 downto 0);
constant int609_t_SLV_LEN : integer := 609;
function int609_t_to_slv(x : int609_t) return std_logic_vector;
function slv_to_int609_t(x : std_logic_vector) return int609_t;
subtype uint610_t is unsigned(609 downto 0);
constant uint610_t_SLV_LEN : integer := 610;
function uint610_t_to_slv(x : uint610_t) return std_logic_vector;
function slv_to_uint610_t(x : std_logic_vector) return uint610_t;
subtype int610_t is signed(609 downto 0);
constant int610_t_SLV_LEN : integer := 610;
function int610_t_to_slv(x : int610_t) return std_logic_vector;
function slv_to_int610_t(x : std_logic_vector) return int610_t;
subtype uint611_t is unsigned(610 downto 0);
constant uint611_t_SLV_LEN : integer := 611;
function uint611_t_to_slv(x : uint611_t) return std_logic_vector;
function slv_to_uint611_t(x : std_logic_vector) return uint611_t;
subtype int611_t is signed(610 downto 0);
constant int611_t_SLV_LEN : integer := 611;
function int611_t_to_slv(x : int611_t) return std_logic_vector;
function slv_to_int611_t(x : std_logic_vector) return int611_t;
subtype uint612_t is unsigned(611 downto 0);
constant uint612_t_SLV_LEN : integer := 612;
function uint612_t_to_slv(x : uint612_t) return std_logic_vector;
function slv_to_uint612_t(x : std_logic_vector) return uint612_t;
subtype int612_t is signed(611 downto 0);
constant int612_t_SLV_LEN : integer := 612;
function int612_t_to_slv(x : int612_t) return std_logic_vector;
function slv_to_int612_t(x : std_logic_vector) return int612_t;
subtype uint613_t is unsigned(612 downto 0);
constant uint613_t_SLV_LEN : integer := 613;
function uint613_t_to_slv(x : uint613_t) return std_logic_vector;
function slv_to_uint613_t(x : std_logic_vector) return uint613_t;
subtype int613_t is signed(612 downto 0);
constant int613_t_SLV_LEN : integer := 613;
function int613_t_to_slv(x : int613_t) return std_logic_vector;
function slv_to_int613_t(x : std_logic_vector) return int613_t;
subtype uint614_t is unsigned(613 downto 0);
constant uint614_t_SLV_LEN : integer := 614;
function uint614_t_to_slv(x : uint614_t) return std_logic_vector;
function slv_to_uint614_t(x : std_logic_vector) return uint614_t;
subtype int614_t is signed(613 downto 0);
constant int614_t_SLV_LEN : integer := 614;
function int614_t_to_slv(x : int614_t) return std_logic_vector;
function slv_to_int614_t(x : std_logic_vector) return int614_t;
subtype uint615_t is unsigned(614 downto 0);
constant uint615_t_SLV_LEN : integer := 615;
function uint615_t_to_slv(x : uint615_t) return std_logic_vector;
function slv_to_uint615_t(x : std_logic_vector) return uint615_t;
subtype int615_t is signed(614 downto 0);
constant int615_t_SLV_LEN : integer := 615;
function int615_t_to_slv(x : int615_t) return std_logic_vector;
function slv_to_int615_t(x : std_logic_vector) return int615_t;
subtype uint616_t is unsigned(615 downto 0);
constant uint616_t_SLV_LEN : integer := 616;
function uint616_t_to_slv(x : uint616_t) return std_logic_vector;
function slv_to_uint616_t(x : std_logic_vector) return uint616_t;
subtype int616_t is signed(615 downto 0);
constant int616_t_SLV_LEN : integer := 616;
function int616_t_to_slv(x : int616_t) return std_logic_vector;
function slv_to_int616_t(x : std_logic_vector) return int616_t;
subtype uint617_t is unsigned(616 downto 0);
constant uint617_t_SLV_LEN : integer := 617;
function uint617_t_to_slv(x : uint617_t) return std_logic_vector;
function slv_to_uint617_t(x : std_logic_vector) return uint617_t;
subtype int617_t is signed(616 downto 0);
constant int617_t_SLV_LEN : integer := 617;
function int617_t_to_slv(x : int617_t) return std_logic_vector;
function slv_to_int617_t(x : std_logic_vector) return int617_t;
subtype uint618_t is unsigned(617 downto 0);
constant uint618_t_SLV_LEN : integer := 618;
function uint618_t_to_slv(x : uint618_t) return std_logic_vector;
function slv_to_uint618_t(x : std_logic_vector) return uint618_t;
subtype int618_t is signed(617 downto 0);
constant int618_t_SLV_LEN : integer := 618;
function int618_t_to_slv(x : int618_t) return std_logic_vector;
function slv_to_int618_t(x : std_logic_vector) return int618_t;
subtype uint619_t is unsigned(618 downto 0);
constant uint619_t_SLV_LEN : integer := 619;
function uint619_t_to_slv(x : uint619_t) return std_logic_vector;
function slv_to_uint619_t(x : std_logic_vector) return uint619_t;
subtype int619_t is signed(618 downto 0);
constant int619_t_SLV_LEN : integer := 619;
function int619_t_to_slv(x : int619_t) return std_logic_vector;
function slv_to_int619_t(x : std_logic_vector) return int619_t;
subtype uint620_t is unsigned(619 downto 0);
constant uint620_t_SLV_LEN : integer := 620;
function uint620_t_to_slv(x : uint620_t) return std_logic_vector;
function slv_to_uint620_t(x : std_logic_vector) return uint620_t;
subtype int620_t is signed(619 downto 0);
constant int620_t_SLV_LEN : integer := 620;
function int620_t_to_slv(x : int620_t) return std_logic_vector;
function slv_to_int620_t(x : std_logic_vector) return int620_t;
subtype uint621_t is unsigned(620 downto 0);
constant uint621_t_SLV_LEN : integer := 621;
function uint621_t_to_slv(x : uint621_t) return std_logic_vector;
function slv_to_uint621_t(x : std_logic_vector) return uint621_t;
subtype int621_t is signed(620 downto 0);
constant int621_t_SLV_LEN : integer := 621;
function int621_t_to_slv(x : int621_t) return std_logic_vector;
function slv_to_int621_t(x : std_logic_vector) return int621_t;
subtype uint622_t is unsigned(621 downto 0);
constant uint622_t_SLV_LEN : integer := 622;
function uint622_t_to_slv(x : uint622_t) return std_logic_vector;
function slv_to_uint622_t(x : std_logic_vector) return uint622_t;
subtype int622_t is signed(621 downto 0);
constant int622_t_SLV_LEN : integer := 622;
function int622_t_to_slv(x : int622_t) return std_logic_vector;
function slv_to_int622_t(x : std_logic_vector) return int622_t;
subtype uint623_t is unsigned(622 downto 0);
constant uint623_t_SLV_LEN : integer := 623;
function uint623_t_to_slv(x : uint623_t) return std_logic_vector;
function slv_to_uint623_t(x : std_logic_vector) return uint623_t;
subtype int623_t is signed(622 downto 0);
constant int623_t_SLV_LEN : integer := 623;
function int623_t_to_slv(x : int623_t) return std_logic_vector;
function slv_to_int623_t(x : std_logic_vector) return int623_t;
subtype uint624_t is unsigned(623 downto 0);
constant uint624_t_SLV_LEN : integer := 624;
function uint624_t_to_slv(x : uint624_t) return std_logic_vector;
function slv_to_uint624_t(x : std_logic_vector) return uint624_t;
subtype int624_t is signed(623 downto 0);
constant int624_t_SLV_LEN : integer := 624;
function int624_t_to_slv(x : int624_t) return std_logic_vector;
function slv_to_int624_t(x : std_logic_vector) return int624_t;
subtype uint625_t is unsigned(624 downto 0);
constant uint625_t_SLV_LEN : integer := 625;
function uint625_t_to_slv(x : uint625_t) return std_logic_vector;
function slv_to_uint625_t(x : std_logic_vector) return uint625_t;
subtype int625_t is signed(624 downto 0);
constant int625_t_SLV_LEN : integer := 625;
function int625_t_to_slv(x : int625_t) return std_logic_vector;
function slv_to_int625_t(x : std_logic_vector) return int625_t;
subtype uint626_t is unsigned(625 downto 0);
constant uint626_t_SLV_LEN : integer := 626;
function uint626_t_to_slv(x : uint626_t) return std_logic_vector;
function slv_to_uint626_t(x : std_logic_vector) return uint626_t;
subtype int626_t is signed(625 downto 0);
constant int626_t_SLV_LEN : integer := 626;
function int626_t_to_slv(x : int626_t) return std_logic_vector;
function slv_to_int626_t(x : std_logic_vector) return int626_t;
subtype uint627_t is unsigned(626 downto 0);
constant uint627_t_SLV_LEN : integer := 627;
function uint627_t_to_slv(x : uint627_t) return std_logic_vector;
function slv_to_uint627_t(x : std_logic_vector) return uint627_t;
subtype int627_t is signed(626 downto 0);
constant int627_t_SLV_LEN : integer := 627;
function int627_t_to_slv(x : int627_t) return std_logic_vector;
function slv_to_int627_t(x : std_logic_vector) return int627_t;
subtype uint628_t is unsigned(627 downto 0);
constant uint628_t_SLV_LEN : integer := 628;
function uint628_t_to_slv(x : uint628_t) return std_logic_vector;
function slv_to_uint628_t(x : std_logic_vector) return uint628_t;
subtype int628_t is signed(627 downto 0);
constant int628_t_SLV_LEN : integer := 628;
function int628_t_to_slv(x : int628_t) return std_logic_vector;
function slv_to_int628_t(x : std_logic_vector) return int628_t;
subtype uint629_t is unsigned(628 downto 0);
constant uint629_t_SLV_LEN : integer := 629;
function uint629_t_to_slv(x : uint629_t) return std_logic_vector;
function slv_to_uint629_t(x : std_logic_vector) return uint629_t;
subtype int629_t is signed(628 downto 0);
constant int629_t_SLV_LEN : integer := 629;
function int629_t_to_slv(x : int629_t) return std_logic_vector;
function slv_to_int629_t(x : std_logic_vector) return int629_t;
subtype uint630_t is unsigned(629 downto 0);
constant uint630_t_SLV_LEN : integer := 630;
function uint630_t_to_slv(x : uint630_t) return std_logic_vector;
function slv_to_uint630_t(x : std_logic_vector) return uint630_t;
subtype int630_t is signed(629 downto 0);
constant int630_t_SLV_LEN : integer := 630;
function int630_t_to_slv(x : int630_t) return std_logic_vector;
function slv_to_int630_t(x : std_logic_vector) return int630_t;
subtype uint631_t is unsigned(630 downto 0);
constant uint631_t_SLV_LEN : integer := 631;
function uint631_t_to_slv(x : uint631_t) return std_logic_vector;
function slv_to_uint631_t(x : std_logic_vector) return uint631_t;
subtype int631_t is signed(630 downto 0);
constant int631_t_SLV_LEN : integer := 631;
function int631_t_to_slv(x : int631_t) return std_logic_vector;
function slv_to_int631_t(x : std_logic_vector) return int631_t;
subtype uint632_t is unsigned(631 downto 0);
constant uint632_t_SLV_LEN : integer := 632;
function uint632_t_to_slv(x : uint632_t) return std_logic_vector;
function slv_to_uint632_t(x : std_logic_vector) return uint632_t;
subtype int632_t is signed(631 downto 0);
constant int632_t_SLV_LEN : integer := 632;
function int632_t_to_slv(x : int632_t) return std_logic_vector;
function slv_to_int632_t(x : std_logic_vector) return int632_t;
subtype uint633_t is unsigned(632 downto 0);
constant uint633_t_SLV_LEN : integer := 633;
function uint633_t_to_slv(x : uint633_t) return std_logic_vector;
function slv_to_uint633_t(x : std_logic_vector) return uint633_t;
subtype int633_t is signed(632 downto 0);
constant int633_t_SLV_LEN : integer := 633;
function int633_t_to_slv(x : int633_t) return std_logic_vector;
function slv_to_int633_t(x : std_logic_vector) return int633_t;
subtype uint634_t is unsigned(633 downto 0);
constant uint634_t_SLV_LEN : integer := 634;
function uint634_t_to_slv(x : uint634_t) return std_logic_vector;
function slv_to_uint634_t(x : std_logic_vector) return uint634_t;
subtype int634_t is signed(633 downto 0);
constant int634_t_SLV_LEN : integer := 634;
function int634_t_to_slv(x : int634_t) return std_logic_vector;
function slv_to_int634_t(x : std_logic_vector) return int634_t;
subtype uint635_t is unsigned(634 downto 0);
constant uint635_t_SLV_LEN : integer := 635;
function uint635_t_to_slv(x : uint635_t) return std_logic_vector;
function slv_to_uint635_t(x : std_logic_vector) return uint635_t;
subtype int635_t is signed(634 downto 0);
constant int635_t_SLV_LEN : integer := 635;
function int635_t_to_slv(x : int635_t) return std_logic_vector;
function slv_to_int635_t(x : std_logic_vector) return int635_t;
subtype uint636_t is unsigned(635 downto 0);
constant uint636_t_SLV_LEN : integer := 636;
function uint636_t_to_slv(x : uint636_t) return std_logic_vector;
function slv_to_uint636_t(x : std_logic_vector) return uint636_t;
subtype int636_t is signed(635 downto 0);
constant int636_t_SLV_LEN : integer := 636;
function int636_t_to_slv(x : int636_t) return std_logic_vector;
function slv_to_int636_t(x : std_logic_vector) return int636_t;
subtype uint637_t is unsigned(636 downto 0);
constant uint637_t_SLV_LEN : integer := 637;
function uint637_t_to_slv(x : uint637_t) return std_logic_vector;
function slv_to_uint637_t(x : std_logic_vector) return uint637_t;
subtype int637_t is signed(636 downto 0);
constant int637_t_SLV_LEN : integer := 637;
function int637_t_to_slv(x : int637_t) return std_logic_vector;
function slv_to_int637_t(x : std_logic_vector) return int637_t;
subtype uint638_t is unsigned(637 downto 0);
constant uint638_t_SLV_LEN : integer := 638;
function uint638_t_to_slv(x : uint638_t) return std_logic_vector;
function slv_to_uint638_t(x : std_logic_vector) return uint638_t;
subtype int638_t is signed(637 downto 0);
constant int638_t_SLV_LEN : integer := 638;
function int638_t_to_slv(x : int638_t) return std_logic_vector;
function slv_to_int638_t(x : std_logic_vector) return int638_t;
subtype uint639_t is unsigned(638 downto 0);
constant uint639_t_SLV_LEN : integer := 639;
function uint639_t_to_slv(x : uint639_t) return std_logic_vector;
function slv_to_uint639_t(x : std_logic_vector) return uint639_t;
subtype int639_t is signed(638 downto 0);
constant int639_t_SLV_LEN : integer := 639;
function int639_t_to_slv(x : int639_t) return std_logic_vector;
function slv_to_int639_t(x : std_logic_vector) return int639_t;
subtype uint640_t is unsigned(639 downto 0);
constant uint640_t_SLV_LEN : integer := 640;
function uint640_t_to_slv(x : uint640_t) return std_logic_vector;
function slv_to_uint640_t(x : std_logic_vector) return uint640_t;
subtype int640_t is signed(639 downto 0);
constant int640_t_SLV_LEN : integer := 640;
function int640_t_to_slv(x : int640_t) return std_logic_vector;
function slv_to_int640_t(x : std_logic_vector) return int640_t;
subtype uint641_t is unsigned(640 downto 0);
constant uint641_t_SLV_LEN : integer := 641;
function uint641_t_to_slv(x : uint641_t) return std_logic_vector;
function slv_to_uint641_t(x : std_logic_vector) return uint641_t;
subtype int641_t is signed(640 downto 0);
constant int641_t_SLV_LEN : integer := 641;
function int641_t_to_slv(x : int641_t) return std_logic_vector;
function slv_to_int641_t(x : std_logic_vector) return int641_t;
subtype uint642_t is unsigned(641 downto 0);
constant uint642_t_SLV_LEN : integer := 642;
function uint642_t_to_slv(x : uint642_t) return std_logic_vector;
function slv_to_uint642_t(x : std_logic_vector) return uint642_t;
subtype int642_t is signed(641 downto 0);
constant int642_t_SLV_LEN : integer := 642;
function int642_t_to_slv(x : int642_t) return std_logic_vector;
function slv_to_int642_t(x : std_logic_vector) return int642_t;
subtype uint643_t is unsigned(642 downto 0);
constant uint643_t_SLV_LEN : integer := 643;
function uint643_t_to_slv(x : uint643_t) return std_logic_vector;
function slv_to_uint643_t(x : std_logic_vector) return uint643_t;
subtype int643_t is signed(642 downto 0);
constant int643_t_SLV_LEN : integer := 643;
function int643_t_to_slv(x : int643_t) return std_logic_vector;
function slv_to_int643_t(x : std_logic_vector) return int643_t;
subtype uint644_t is unsigned(643 downto 0);
constant uint644_t_SLV_LEN : integer := 644;
function uint644_t_to_slv(x : uint644_t) return std_logic_vector;
function slv_to_uint644_t(x : std_logic_vector) return uint644_t;
subtype int644_t is signed(643 downto 0);
constant int644_t_SLV_LEN : integer := 644;
function int644_t_to_slv(x : int644_t) return std_logic_vector;
function slv_to_int644_t(x : std_logic_vector) return int644_t;
subtype uint645_t is unsigned(644 downto 0);
constant uint645_t_SLV_LEN : integer := 645;
function uint645_t_to_slv(x : uint645_t) return std_logic_vector;
function slv_to_uint645_t(x : std_logic_vector) return uint645_t;
subtype int645_t is signed(644 downto 0);
constant int645_t_SLV_LEN : integer := 645;
function int645_t_to_slv(x : int645_t) return std_logic_vector;
function slv_to_int645_t(x : std_logic_vector) return int645_t;
subtype uint646_t is unsigned(645 downto 0);
constant uint646_t_SLV_LEN : integer := 646;
function uint646_t_to_slv(x : uint646_t) return std_logic_vector;
function slv_to_uint646_t(x : std_logic_vector) return uint646_t;
subtype int646_t is signed(645 downto 0);
constant int646_t_SLV_LEN : integer := 646;
function int646_t_to_slv(x : int646_t) return std_logic_vector;
function slv_to_int646_t(x : std_logic_vector) return int646_t;
subtype uint647_t is unsigned(646 downto 0);
constant uint647_t_SLV_LEN : integer := 647;
function uint647_t_to_slv(x : uint647_t) return std_logic_vector;
function slv_to_uint647_t(x : std_logic_vector) return uint647_t;
subtype int647_t is signed(646 downto 0);
constant int647_t_SLV_LEN : integer := 647;
function int647_t_to_slv(x : int647_t) return std_logic_vector;
function slv_to_int647_t(x : std_logic_vector) return int647_t;
subtype uint648_t is unsigned(647 downto 0);
constant uint648_t_SLV_LEN : integer := 648;
function uint648_t_to_slv(x : uint648_t) return std_logic_vector;
function slv_to_uint648_t(x : std_logic_vector) return uint648_t;
subtype int648_t is signed(647 downto 0);
constant int648_t_SLV_LEN : integer := 648;
function int648_t_to_slv(x : int648_t) return std_logic_vector;
function slv_to_int648_t(x : std_logic_vector) return int648_t;
subtype uint649_t is unsigned(648 downto 0);
constant uint649_t_SLV_LEN : integer := 649;
function uint649_t_to_slv(x : uint649_t) return std_logic_vector;
function slv_to_uint649_t(x : std_logic_vector) return uint649_t;
subtype int649_t is signed(648 downto 0);
constant int649_t_SLV_LEN : integer := 649;
function int649_t_to_slv(x : int649_t) return std_logic_vector;
function slv_to_int649_t(x : std_logic_vector) return int649_t;
subtype uint650_t is unsigned(649 downto 0);
constant uint650_t_SLV_LEN : integer := 650;
function uint650_t_to_slv(x : uint650_t) return std_logic_vector;
function slv_to_uint650_t(x : std_logic_vector) return uint650_t;
subtype int650_t is signed(649 downto 0);
constant int650_t_SLV_LEN : integer := 650;
function int650_t_to_slv(x : int650_t) return std_logic_vector;
function slv_to_int650_t(x : std_logic_vector) return int650_t;
subtype uint651_t is unsigned(650 downto 0);
constant uint651_t_SLV_LEN : integer := 651;
function uint651_t_to_slv(x : uint651_t) return std_logic_vector;
function slv_to_uint651_t(x : std_logic_vector) return uint651_t;
subtype int651_t is signed(650 downto 0);
constant int651_t_SLV_LEN : integer := 651;
function int651_t_to_slv(x : int651_t) return std_logic_vector;
function slv_to_int651_t(x : std_logic_vector) return int651_t;
subtype uint652_t is unsigned(651 downto 0);
constant uint652_t_SLV_LEN : integer := 652;
function uint652_t_to_slv(x : uint652_t) return std_logic_vector;
function slv_to_uint652_t(x : std_logic_vector) return uint652_t;
subtype int652_t is signed(651 downto 0);
constant int652_t_SLV_LEN : integer := 652;
function int652_t_to_slv(x : int652_t) return std_logic_vector;
function slv_to_int652_t(x : std_logic_vector) return int652_t;
subtype uint653_t is unsigned(652 downto 0);
constant uint653_t_SLV_LEN : integer := 653;
function uint653_t_to_slv(x : uint653_t) return std_logic_vector;
function slv_to_uint653_t(x : std_logic_vector) return uint653_t;
subtype int653_t is signed(652 downto 0);
constant int653_t_SLV_LEN : integer := 653;
function int653_t_to_slv(x : int653_t) return std_logic_vector;
function slv_to_int653_t(x : std_logic_vector) return int653_t;
subtype uint654_t is unsigned(653 downto 0);
constant uint654_t_SLV_LEN : integer := 654;
function uint654_t_to_slv(x : uint654_t) return std_logic_vector;
function slv_to_uint654_t(x : std_logic_vector) return uint654_t;
subtype int654_t is signed(653 downto 0);
constant int654_t_SLV_LEN : integer := 654;
function int654_t_to_slv(x : int654_t) return std_logic_vector;
function slv_to_int654_t(x : std_logic_vector) return int654_t;
subtype uint655_t is unsigned(654 downto 0);
constant uint655_t_SLV_LEN : integer := 655;
function uint655_t_to_slv(x : uint655_t) return std_logic_vector;
function slv_to_uint655_t(x : std_logic_vector) return uint655_t;
subtype int655_t is signed(654 downto 0);
constant int655_t_SLV_LEN : integer := 655;
function int655_t_to_slv(x : int655_t) return std_logic_vector;
function slv_to_int655_t(x : std_logic_vector) return int655_t;
subtype uint656_t is unsigned(655 downto 0);
constant uint656_t_SLV_LEN : integer := 656;
function uint656_t_to_slv(x : uint656_t) return std_logic_vector;
function slv_to_uint656_t(x : std_logic_vector) return uint656_t;
subtype int656_t is signed(655 downto 0);
constant int656_t_SLV_LEN : integer := 656;
function int656_t_to_slv(x : int656_t) return std_logic_vector;
function slv_to_int656_t(x : std_logic_vector) return int656_t;
subtype uint657_t is unsigned(656 downto 0);
constant uint657_t_SLV_LEN : integer := 657;
function uint657_t_to_slv(x : uint657_t) return std_logic_vector;
function slv_to_uint657_t(x : std_logic_vector) return uint657_t;
subtype int657_t is signed(656 downto 0);
constant int657_t_SLV_LEN : integer := 657;
function int657_t_to_slv(x : int657_t) return std_logic_vector;
function slv_to_int657_t(x : std_logic_vector) return int657_t;
subtype uint658_t is unsigned(657 downto 0);
constant uint658_t_SLV_LEN : integer := 658;
function uint658_t_to_slv(x : uint658_t) return std_logic_vector;
function slv_to_uint658_t(x : std_logic_vector) return uint658_t;
subtype int658_t is signed(657 downto 0);
constant int658_t_SLV_LEN : integer := 658;
function int658_t_to_slv(x : int658_t) return std_logic_vector;
function slv_to_int658_t(x : std_logic_vector) return int658_t;
subtype uint659_t is unsigned(658 downto 0);
constant uint659_t_SLV_LEN : integer := 659;
function uint659_t_to_slv(x : uint659_t) return std_logic_vector;
function slv_to_uint659_t(x : std_logic_vector) return uint659_t;
subtype int659_t is signed(658 downto 0);
constant int659_t_SLV_LEN : integer := 659;
function int659_t_to_slv(x : int659_t) return std_logic_vector;
function slv_to_int659_t(x : std_logic_vector) return int659_t;
subtype uint660_t is unsigned(659 downto 0);
constant uint660_t_SLV_LEN : integer := 660;
function uint660_t_to_slv(x : uint660_t) return std_logic_vector;
function slv_to_uint660_t(x : std_logic_vector) return uint660_t;
subtype int660_t is signed(659 downto 0);
constant int660_t_SLV_LEN : integer := 660;
function int660_t_to_slv(x : int660_t) return std_logic_vector;
function slv_to_int660_t(x : std_logic_vector) return int660_t;
subtype uint661_t is unsigned(660 downto 0);
constant uint661_t_SLV_LEN : integer := 661;
function uint661_t_to_slv(x : uint661_t) return std_logic_vector;
function slv_to_uint661_t(x : std_logic_vector) return uint661_t;
subtype int661_t is signed(660 downto 0);
constant int661_t_SLV_LEN : integer := 661;
function int661_t_to_slv(x : int661_t) return std_logic_vector;
function slv_to_int661_t(x : std_logic_vector) return int661_t;
subtype uint662_t is unsigned(661 downto 0);
constant uint662_t_SLV_LEN : integer := 662;
function uint662_t_to_slv(x : uint662_t) return std_logic_vector;
function slv_to_uint662_t(x : std_logic_vector) return uint662_t;
subtype int662_t is signed(661 downto 0);
constant int662_t_SLV_LEN : integer := 662;
function int662_t_to_slv(x : int662_t) return std_logic_vector;
function slv_to_int662_t(x : std_logic_vector) return int662_t;
subtype uint663_t is unsigned(662 downto 0);
constant uint663_t_SLV_LEN : integer := 663;
function uint663_t_to_slv(x : uint663_t) return std_logic_vector;
function slv_to_uint663_t(x : std_logic_vector) return uint663_t;
subtype int663_t is signed(662 downto 0);
constant int663_t_SLV_LEN : integer := 663;
function int663_t_to_slv(x : int663_t) return std_logic_vector;
function slv_to_int663_t(x : std_logic_vector) return int663_t;
subtype uint664_t is unsigned(663 downto 0);
constant uint664_t_SLV_LEN : integer := 664;
function uint664_t_to_slv(x : uint664_t) return std_logic_vector;
function slv_to_uint664_t(x : std_logic_vector) return uint664_t;
subtype int664_t is signed(663 downto 0);
constant int664_t_SLV_LEN : integer := 664;
function int664_t_to_slv(x : int664_t) return std_logic_vector;
function slv_to_int664_t(x : std_logic_vector) return int664_t;
subtype uint665_t is unsigned(664 downto 0);
constant uint665_t_SLV_LEN : integer := 665;
function uint665_t_to_slv(x : uint665_t) return std_logic_vector;
function slv_to_uint665_t(x : std_logic_vector) return uint665_t;
subtype int665_t is signed(664 downto 0);
constant int665_t_SLV_LEN : integer := 665;
function int665_t_to_slv(x : int665_t) return std_logic_vector;
function slv_to_int665_t(x : std_logic_vector) return int665_t;
subtype uint666_t is unsigned(665 downto 0);
constant uint666_t_SLV_LEN : integer := 666;
function uint666_t_to_slv(x : uint666_t) return std_logic_vector;
function slv_to_uint666_t(x : std_logic_vector) return uint666_t;
subtype int666_t is signed(665 downto 0);
constant int666_t_SLV_LEN : integer := 666;
function int666_t_to_slv(x : int666_t) return std_logic_vector;
function slv_to_int666_t(x : std_logic_vector) return int666_t;
subtype uint667_t is unsigned(666 downto 0);
constant uint667_t_SLV_LEN : integer := 667;
function uint667_t_to_slv(x : uint667_t) return std_logic_vector;
function slv_to_uint667_t(x : std_logic_vector) return uint667_t;
subtype int667_t is signed(666 downto 0);
constant int667_t_SLV_LEN : integer := 667;
function int667_t_to_slv(x : int667_t) return std_logic_vector;
function slv_to_int667_t(x : std_logic_vector) return int667_t;
subtype uint668_t is unsigned(667 downto 0);
constant uint668_t_SLV_LEN : integer := 668;
function uint668_t_to_slv(x : uint668_t) return std_logic_vector;
function slv_to_uint668_t(x : std_logic_vector) return uint668_t;
subtype int668_t is signed(667 downto 0);
constant int668_t_SLV_LEN : integer := 668;
function int668_t_to_slv(x : int668_t) return std_logic_vector;
function slv_to_int668_t(x : std_logic_vector) return int668_t;
subtype uint669_t is unsigned(668 downto 0);
constant uint669_t_SLV_LEN : integer := 669;
function uint669_t_to_slv(x : uint669_t) return std_logic_vector;
function slv_to_uint669_t(x : std_logic_vector) return uint669_t;
subtype int669_t is signed(668 downto 0);
constant int669_t_SLV_LEN : integer := 669;
function int669_t_to_slv(x : int669_t) return std_logic_vector;
function slv_to_int669_t(x : std_logic_vector) return int669_t;
subtype uint670_t is unsigned(669 downto 0);
constant uint670_t_SLV_LEN : integer := 670;
function uint670_t_to_slv(x : uint670_t) return std_logic_vector;
function slv_to_uint670_t(x : std_logic_vector) return uint670_t;
subtype int670_t is signed(669 downto 0);
constant int670_t_SLV_LEN : integer := 670;
function int670_t_to_slv(x : int670_t) return std_logic_vector;
function slv_to_int670_t(x : std_logic_vector) return int670_t;
subtype uint671_t is unsigned(670 downto 0);
constant uint671_t_SLV_LEN : integer := 671;
function uint671_t_to_slv(x : uint671_t) return std_logic_vector;
function slv_to_uint671_t(x : std_logic_vector) return uint671_t;
subtype int671_t is signed(670 downto 0);
constant int671_t_SLV_LEN : integer := 671;
function int671_t_to_slv(x : int671_t) return std_logic_vector;
function slv_to_int671_t(x : std_logic_vector) return int671_t;
subtype uint672_t is unsigned(671 downto 0);
constant uint672_t_SLV_LEN : integer := 672;
function uint672_t_to_slv(x : uint672_t) return std_logic_vector;
function slv_to_uint672_t(x : std_logic_vector) return uint672_t;
subtype int672_t is signed(671 downto 0);
constant int672_t_SLV_LEN : integer := 672;
function int672_t_to_slv(x : int672_t) return std_logic_vector;
function slv_to_int672_t(x : std_logic_vector) return int672_t;
subtype uint673_t is unsigned(672 downto 0);
constant uint673_t_SLV_LEN : integer := 673;
function uint673_t_to_slv(x : uint673_t) return std_logic_vector;
function slv_to_uint673_t(x : std_logic_vector) return uint673_t;
subtype int673_t is signed(672 downto 0);
constant int673_t_SLV_LEN : integer := 673;
function int673_t_to_slv(x : int673_t) return std_logic_vector;
function slv_to_int673_t(x : std_logic_vector) return int673_t;
subtype uint674_t is unsigned(673 downto 0);
constant uint674_t_SLV_LEN : integer := 674;
function uint674_t_to_slv(x : uint674_t) return std_logic_vector;
function slv_to_uint674_t(x : std_logic_vector) return uint674_t;
subtype int674_t is signed(673 downto 0);
constant int674_t_SLV_LEN : integer := 674;
function int674_t_to_slv(x : int674_t) return std_logic_vector;
function slv_to_int674_t(x : std_logic_vector) return int674_t;
subtype uint675_t is unsigned(674 downto 0);
constant uint675_t_SLV_LEN : integer := 675;
function uint675_t_to_slv(x : uint675_t) return std_logic_vector;
function slv_to_uint675_t(x : std_logic_vector) return uint675_t;
subtype int675_t is signed(674 downto 0);
constant int675_t_SLV_LEN : integer := 675;
function int675_t_to_slv(x : int675_t) return std_logic_vector;
function slv_to_int675_t(x : std_logic_vector) return int675_t;
subtype uint676_t is unsigned(675 downto 0);
constant uint676_t_SLV_LEN : integer := 676;
function uint676_t_to_slv(x : uint676_t) return std_logic_vector;
function slv_to_uint676_t(x : std_logic_vector) return uint676_t;
subtype int676_t is signed(675 downto 0);
constant int676_t_SLV_LEN : integer := 676;
function int676_t_to_slv(x : int676_t) return std_logic_vector;
function slv_to_int676_t(x : std_logic_vector) return int676_t;
subtype uint677_t is unsigned(676 downto 0);
constant uint677_t_SLV_LEN : integer := 677;
function uint677_t_to_slv(x : uint677_t) return std_logic_vector;
function slv_to_uint677_t(x : std_logic_vector) return uint677_t;
subtype int677_t is signed(676 downto 0);
constant int677_t_SLV_LEN : integer := 677;
function int677_t_to_slv(x : int677_t) return std_logic_vector;
function slv_to_int677_t(x : std_logic_vector) return int677_t;
subtype uint678_t is unsigned(677 downto 0);
constant uint678_t_SLV_LEN : integer := 678;
function uint678_t_to_slv(x : uint678_t) return std_logic_vector;
function slv_to_uint678_t(x : std_logic_vector) return uint678_t;
subtype int678_t is signed(677 downto 0);
constant int678_t_SLV_LEN : integer := 678;
function int678_t_to_slv(x : int678_t) return std_logic_vector;
function slv_to_int678_t(x : std_logic_vector) return int678_t;
subtype uint679_t is unsigned(678 downto 0);
constant uint679_t_SLV_LEN : integer := 679;
function uint679_t_to_slv(x : uint679_t) return std_logic_vector;
function slv_to_uint679_t(x : std_logic_vector) return uint679_t;
subtype int679_t is signed(678 downto 0);
constant int679_t_SLV_LEN : integer := 679;
function int679_t_to_slv(x : int679_t) return std_logic_vector;
function slv_to_int679_t(x : std_logic_vector) return int679_t;
subtype uint680_t is unsigned(679 downto 0);
constant uint680_t_SLV_LEN : integer := 680;
function uint680_t_to_slv(x : uint680_t) return std_logic_vector;
function slv_to_uint680_t(x : std_logic_vector) return uint680_t;
subtype int680_t is signed(679 downto 0);
constant int680_t_SLV_LEN : integer := 680;
function int680_t_to_slv(x : int680_t) return std_logic_vector;
function slv_to_int680_t(x : std_logic_vector) return int680_t;
subtype uint681_t is unsigned(680 downto 0);
constant uint681_t_SLV_LEN : integer := 681;
function uint681_t_to_slv(x : uint681_t) return std_logic_vector;
function slv_to_uint681_t(x : std_logic_vector) return uint681_t;
subtype int681_t is signed(680 downto 0);
constant int681_t_SLV_LEN : integer := 681;
function int681_t_to_slv(x : int681_t) return std_logic_vector;
function slv_to_int681_t(x : std_logic_vector) return int681_t;
subtype uint682_t is unsigned(681 downto 0);
constant uint682_t_SLV_LEN : integer := 682;
function uint682_t_to_slv(x : uint682_t) return std_logic_vector;
function slv_to_uint682_t(x : std_logic_vector) return uint682_t;
subtype int682_t is signed(681 downto 0);
constant int682_t_SLV_LEN : integer := 682;
function int682_t_to_slv(x : int682_t) return std_logic_vector;
function slv_to_int682_t(x : std_logic_vector) return int682_t;
subtype uint683_t is unsigned(682 downto 0);
constant uint683_t_SLV_LEN : integer := 683;
function uint683_t_to_slv(x : uint683_t) return std_logic_vector;
function slv_to_uint683_t(x : std_logic_vector) return uint683_t;
subtype int683_t is signed(682 downto 0);
constant int683_t_SLV_LEN : integer := 683;
function int683_t_to_slv(x : int683_t) return std_logic_vector;
function slv_to_int683_t(x : std_logic_vector) return int683_t;
subtype uint684_t is unsigned(683 downto 0);
constant uint684_t_SLV_LEN : integer := 684;
function uint684_t_to_slv(x : uint684_t) return std_logic_vector;
function slv_to_uint684_t(x : std_logic_vector) return uint684_t;
subtype int684_t is signed(683 downto 0);
constant int684_t_SLV_LEN : integer := 684;
function int684_t_to_slv(x : int684_t) return std_logic_vector;
function slv_to_int684_t(x : std_logic_vector) return int684_t;
subtype uint685_t is unsigned(684 downto 0);
constant uint685_t_SLV_LEN : integer := 685;
function uint685_t_to_slv(x : uint685_t) return std_logic_vector;
function slv_to_uint685_t(x : std_logic_vector) return uint685_t;
subtype int685_t is signed(684 downto 0);
constant int685_t_SLV_LEN : integer := 685;
function int685_t_to_slv(x : int685_t) return std_logic_vector;
function slv_to_int685_t(x : std_logic_vector) return int685_t;
subtype uint686_t is unsigned(685 downto 0);
constant uint686_t_SLV_LEN : integer := 686;
function uint686_t_to_slv(x : uint686_t) return std_logic_vector;
function slv_to_uint686_t(x : std_logic_vector) return uint686_t;
subtype int686_t is signed(685 downto 0);
constant int686_t_SLV_LEN : integer := 686;
function int686_t_to_slv(x : int686_t) return std_logic_vector;
function slv_to_int686_t(x : std_logic_vector) return int686_t;
subtype uint687_t is unsigned(686 downto 0);
constant uint687_t_SLV_LEN : integer := 687;
function uint687_t_to_slv(x : uint687_t) return std_logic_vector;
function slv_to_uint687_t(x : std_logic_vector) return uint687_t;
subtype int687_t is signed(686 downto 0);
constant int687_t_SLV_LEN : integer := 687;
function int687_t_to_slv(x : int687_t) return std_logic_vector;
function slv_to_int687_t(x : std_logic_vector) return int687_t;
subtype uint688_t is unsigned(687 downto 0);
constant uint688_t_SLV_LEN : integer := 688;
function uint688_t_to_slv(x : uint688_t) return std_logic_vector;
function slv_to_uint688_t(x : std_logic_vector) return uint688_t;
subtype int688_t is signed(687 downto 0);
constant int688_t_SLV_LEN : integer := 688;
function int688_t_to_slv(x : int688_t) return std_logic_vector;
function slv_to_int688_t(x : std_logic_vector) return int688_t;
subtype uint689_t is unsigned(688 downto 0);
constant uint689_t_SLV_LEN : integer := 689;
function uint689_t_to_slv(x : uint689_t) return std_logic_vector;
function slv_to_uint689_t(x : std_logic_vector) return uint689_t;
subtype int689_t is signed(688 downto 0);
constant int689_t_SLV_LEN : integer := 689;
function int689_t_to_slv(x : int689_t) return std_logic_vector;
function slv_to_int689_t(x : std_logic_vector) return int689_t;
subtype uint690_t is unsigned(689 downto 0);
constant uint690_t_SLV_LEN : integer := 690;
function uint690_t_to_slv(x : uint690_t) return std_logic_vector;
function slv_to_uint690_t(x : std_logic_vector) return uint690_t;
subtype int690_t is signed(689 downto 0);
constant int690_t_SLV_LEN : integer := 690;
function int690_t_to_slv(x : int690_t) return std_logic_vector;
function slv_to_int690_t(x : std_logic_vector) return int690_t;
subtype uint691_t is unsigned(690 downto 0);
constant uint691_t_SLV_LEN : integer := 691;
function uint691_t_to_slv(x : uint691_t) return std_logic_vector;
function slv_to_uint691_t(x : std_logic_vector) return uint691_t;
subtype int691_t is signed(690 downto 0);
constant int691_t_SLV_LEN : integer := 691;
function int691_t_to_slv(x : int691_t) return std_logic_vector;
function slv_to_int691_t(x : std_logic_vector) return int691_t;
subtype uint692_t is unsigned(691 downto 0);
constant uint692_t_SLV_LEN : integer := 692;
function uint692_t_to_slv(x : uint692_t) return std_logic_vector;
function slv_to_uint692_t(x : std_logic_vector) return uint692_t;
subtype int692_t is signed(691 downto 0);
constant int692_t_SLV_LEN : integer := 692;
function int692_t_to_slv(x : int692_t) return std_logic_vector;
function slv_to_int692_t(x : std_logic_vector) return int692_t;
subtype uint693_t is unsigned(692 downto 0);
constant uint693_t_SLV_LEN : integer := 693;
function uint693_t_to_slv(x : uint693_t) return std_logic_vector;
function slv_to_uint693_t(x : std_logic_vector) return uint693_t;
subtype int693_t is signed(692 downto 0);
constant int693_t_SLV_LEN : integer := 693;
function int693_t_to_slv(x : int693_t) return std_logic_vector;
function slv_to_int693_t(x : std_logic_vector) return int693_t;
subtype uint694_t is unsigned(693 downto 0);
constant uint694_t_SLV_LEN : integer := 694;
function uint694_t_to_slv(x : uint694_t) return std_logic_vector;
function slv_to_uint694_t(x : std_logic_vector) return uint694_t;
subtype int694_t is signed(693 downto 0);
constant int694_t_SLV_LEN : integer := 694;
function int694_t_to_slv(x : int694_t) return std_logic_vector;
function slv_to_int694_t(x : std_logic_vector) return int694_t;
subtype uint695_t is unsigned(694 downto 0);
constant uint695_t_SLV_LEN : integer := 695;
function uint695_t_to_slv(x : uint695_t) return std_logic_vector;
function slv_to_uint695_t(x : std_logic_vector) return uint695_t;
subtype int695_t is signed(694 downto 0);
constant int695_t_SLV_LEN : integer := 695;
function int695_t_to_slv(x : int695_t) return std_logic_vector;
function slv_to_int695_t(x : std_logic_vector) return int695_t;
subtype uint696_t is unsigned(695 downto 0);
constant uint696_t_SLV_LEN : integer := 696;
function uint696_t_to_slv(x : uint696_t) return std_logic_vector;
function slv_to_uint696_t(x : std_logic_vector) return uint696_t;
subtype int696_t is signed(695 downto 0);
constant int696_t_SLV_LEN : integer := 696;
function int696_t_to_slv(x : int696_t) return std_logic_vector;
function slv_to_int696_t(x : std_logic_vector) return int696_t;
subtype uint697_t is unsigned(696 downto 0);
constant uint697_t_SLV_LEN : integer := 697;
function uint697_t_to_slv(x : uint697_t) return std_logic_vector;
function slv_to_uint697_t(x : std_logic_vector) return uint697_t;
subtype int697_t is signed(696 downto 0);
constant int697_t_SLV_LEN : integer := 697;
function int697_t_to_slv(x : int697_t) return std_logic_vector;
function slv_to_int697_t(x : std_logic_vector) return int697_t;
subtype uint698_t is unsigned(697 downto 0);
constant uint698_t_SLV_LEN : integer := 698;
function uint698_t_to_slv(x : uint698_t) return std_logic_vector;
function slv_to_uint698_t(x : std_logic_vector) return uint698_t;
subtype int698_t is signed(697 downto 0);
constant int698_t_SLV_LEN : integer := 698;
function int698_t_to_slv(x : int698_t) return std_logic_vector;
function slv_to_int698_t(x : std_logic_vector) return int698_t;
subtype uint699_t is unsigned(698 downto 0);
constant uint699_t_SLV_LEN : integer := 699;
function uint699_t_to_slv(x : uint699_t) return std_logic_vector;
function slv_to_uint699_t(x : std_logic_vector) return uint699_t;
subtype int699_t is signed(698 downto 0);
constant int699_t_SLV_LEN : integer := 699;
function int699_t_to_slv(x : int699_t) return std_logic_vector;
function slv_to_int699_t(x : std_logic_vector) return int699_t;
subtype uint700_t is unsigned(699 downto 0);
constant uint700_t_SLV_LEN : integer := 700;
function uint700_t_to_slv(x : uint700_t) return std_logic_vector;
function slv_to_uint700_t(x : std_logic_vector) return uint700_t;
subtype int700_t is signed(699 downto 0);
constant int700_t_SLV_LEN : integer := 700;
function int700_t_to_slv(x : int700_t) return std_logic_vector;
function slv_to_int700_t(x : std_logic_vector) return int700_t;
subtype uint701_t is unsigned(700 downto 0);
constant uint701_t_SLV_LEN : integer := 701;
function uint701_t_to_slv(x : uint701_t) return std_logic_vector;
function slv_to_uint701_t(x : std_logic_vector) return uint701_t;
subtype int701_t is signed(700 downto 0);
constant int701_t_SLV_LEN : integer := 701;
function int701_t_to_slv(x : int701_t) return std_logic_vector;
function slv_to_int701_t(x : std_logic_vector) return int701_t;
subtype uint702_t is unsigned(701 downto 0);
constant uint702_t_SLV_LEN : integer := 702;
function uint702_t_to_slv(x : uint702_t) return std_logic_vector;
function slv_to_uint702_t(x : std_logic_vector) return uint702_t;
subtype int702_t is signed(701 downto 0);
constant int702_t_SLV_LEN : integer := 702;
function int702_t_to_slv(x : int702_t) return std_logic_vector;
function slv_to_int702_t(x : std_logic_vector) return int702_t;
subtype uint703_t is unsigned(702 downto 0);
constant uint703_t_SLV_LEN : integer := 703;
function uint703_t_to_slv(x : uint703_t) return std_logic_vector;
function slv_to_uint703_t(x : std_logic_vector) return uint703_t;
subtype int703_t is signed(702 downto 0);
constant int703_t_SLV_LEN : integer := 703;
function int703_t_to_slv(x : int703_t) return std_logic_vector;
function slv_to_int703_t(x : std_logic_vector) return int703_t;
subtype uint704_t is unsigned(703 downto 0);
constant uint704_t_SLV_LEN : integer := 704;
function uint704_t_to_slv(x : uint704_t) return std_logic_vector;
function slv_to_uint704_t(x : std_logic_vector) return uint704_t;
subtype int704_t is signed(703 downto 0);
constant int704_t_SLV_LEN : integer := 704;
function int704_t_to_slv(x : int704_t) return std_logic_vector;
function slv_to_int704_t(x : std_logic_vector) return int704_t;
subtype uint705_t is unsigned(704 downto 0);
constant uint705_t_SLV_LEN : integer := 705;
function uint705_t_to_slv(x : uint705_t) return std_logic_vector;
function slv_to_uint705_t(x : std_logic_vector) return uint705_t;
subtype int705_t is signed(704 downto 0);
constant int705_t_SLV_LEN : integer := 705;
function int705_t_to_slv(x : int705_t) return std_logic_vector;
function slv_to_int705_t(x : std_logic_vector) return int705_t;
subtype uint706_t is unsigned(705 downto 0);
constant uint706_t_SLV_LEN : integer := 706;
function uint706_t_to_slv(x : uint706_t) return std_logic_vector;
function slv_to_uint706_t(x : std_logic_vector) return uint706_t;
subtype int706_t is signed(705 downto 0);
constant int706_t_SLV_LEN : integer := 706;
function int706_t_to_slv(x : int706_t) return std_logic_vector;
function slv_to_int706_t(x : std_logic_vector) return int706_t;
subtype uint707_t is unsigned(706 downto 0);
constant uint707_t_SLV_LEN : integer := 707;
function uint707_t_to_slv(x : uint707_t) return std_logic_vector;
function slv_to_uint707_t(x : std_logic_vector) return uint707_t;
subtype int707_t is signed(706 downto 0);
constant int707_t_SLV_LEN : integer := 707;
function int707_t_to_slv(x : int707_t) return std_logic_vector;
function slv_to_int707_t(x : std_logic_vector) return int707_t;
subtype uint708_t is unsigned(707 downto 0);
constant uint708_t_SLV_LEN : integer := 708;
function uint708_t_to_slv(x : uint708_t) return std_logic_vector;
function slv_to_uint708_t(x : std_logic_vector) return uint708_t;
subtype int708_t is signed(707 downto 0);
constant int708_t_SLV_LEN : integer := 708;
function int708_t_to_slv(x : int708_t) return std_logic_vector;
function slv_to_int708_t(x : std_logic_vector) return int708_t;
subtype uint709_t is unsigned(708 downto 0);
constant uint709_t_SLV_LEN : integer := 709;
function uint709_t_to_slv(x : uint709_t) return std_logic_vector;
function slv_to_uint709_t(x : std_logic_vector) return uint709_t;
subtype int709_t is signed(708 downto 0);
constant int709_t_SLV_LEN : integer := 709;
function int709_t_to_slv(x : int709_t) return std_logic_vector;
function slv_to_int709_t(x : std_logic_vector) return int709_t;
subtype uint710_t is unsigned(709 downto 0);
constant uint710_t_SLV_LEN : integer := 710;
function uint710_t_to_slv(x : uint710_t) return std_logic_vector;
function slv_to_uint710_t(x : std_logic_vector) return uint710_t;
subtype int710_t is signed(709 downto 0);
constant int710_t_SLV_LEN : integer := 710;
function int710_t_to_slv(x : int710_t) return std_logic_vector;
function slv_to_int710_t(x : std_logic_vector) return int710_t;
subtype uint711_t is unsigned(710 downto 0);
constant uint711_t_SLV_LEN : integer := 711;
function uint711_t_to_slv(x : uint711_t) return std_logic_vector;
function slv_to_uint711_t(x : std_logic_vector) return uint711_t;
subtype int711_t is signed(710 downto 0);
constant int711_t_SLV_LEN : integer := 711;
function int711_t_to_slv(x : int711_t) return std_logic_vector;
function slv_to_int711_t(x : std_logic_vector) return int711_t;
subtype uint712_t is unsigned(711 downto 0);
constant uint712_t_SLV_LEN : integer := 712;
function uint712_t_to_slv(x : uint712_t) return std_logic_vector;
function slv_to_uint712_t(x : std_logic_vector) return uint712_t;
subtype int712_t is signed(711 downto 0);
constant int712_t_SLV_LEN : integer := 712;
function int712_t_to_slv(x : int712_t) return std_logic_vector;
function slv_to_int712_t(x : std_logic_vector) return int712_t;
subtype uint713_t is unsigned(712 downto 0);
constant uint713_t_SLV_LEN : integer := 713;
function uint713_t_to_slv(x : uint713_t) return std_logic_vector;
function slv_to_uint713_t(x : std_logic_vector) return uint713_t;
subtype int713_t is signed(712 downto 0);
constant int713_t_SLV_LEN : integer := 713;
function int713_t_to_slv(x : int713_t) return std_logic_vector;
function slv_to_int713_t(x : std_logic_vector) return int713_t;
subtype uint714_t is unsigned(713 downto 0);
constant uint714_t_SLV_LEN : integer := 714;
function uint714_t_to_slv(x : uint714_t) return std_logic_vector;
function slv_to_uint714_t(x : std_logic_vector) return uint714_t;
subtype int714_t is signed(713 downto 0);
constant int714_t_SLV_LEN : integer := 714;
function int714_t_to_slv(x : int714_t) return std_logic_vector;
function slv_to_int714_t(x : std_logic_vector) return int714_t;
subtype uint715_t is unsigned(714 downto 0);
constant uint715_t_SLV_LEN : integer := 715;
function uint715_t_to_slv(x : uint715_t) return std_logic_vector;
function slv_to_uint715_t(x : std_logic_vector) return uint715_t;
subtype int715_t is signed(714 downto 0);
constant int715_t_SLV_LEN : integer := 715;
function int715_t_to_slv(x : int715_t) return std_logic_vector;
function slv_to_int715_t(x : std_logic_vector) return int715_t;
subtype uint716_t is unsigned(715 downto 0);
constant uint716_t_SLV_LEN : integer := 716;
function uint716_t_to_slv(x : uint716_t) return std_logic_vector;
function slv_to_uint716_t(x : std_logic_vector) return uint716_t;
subtype int716_t is signed(715 downto 0);
constant int716_t_SLV_LEN : integer := 716;
function int716_t_to_slv(x : int716_t) return std_logic_vector;
function slv_to_int716_t(x : std_logic_vector) return int716_t;
subtype uint717_t is unsigned(716 downto 0);
constant uint717_t_SLV_LEN : integer := 717;
function uint717_t_to_slv(x : uint717_t) return std_logic_vector;
function slv_to_uint717_t(x : std_logic_vector) return uint717_t;
subtype int717_t is signed(716 downto 0);
constant int717_t_SLV_LEN : integer := 717;
function int717_t_to_slv(x : int717_t) return std_logic_vector;
function slv_to_int717_t(x : std_logic_vector) return int717_t;
subtype uint718_t is unsigned(717 downto 0);
constant uint718_t_SLV_LEN : integer := 718;
function uint718_t_to_slv(x : uint718_t) return std_logic_vector;
function slv_to_uint718_t(x : std_logic_vector) return uint718_t;
subtype int718_t is signed(717 downto 0);
constant int718_t_SLV_LEN : integer := 718;
function int718_t_to_slv(x : int718_t) return std_logic_vector;
function slv_to_int718_t(x : std_logic_vector) return int718_t;
subtype uint719_t is unsigned(718 downto 0);
constant uint719_t_SLV_LEN : integer := 719;
function uint719_t_to_slv(x : uint719_t) return std_logic_vector;
function slv_to_uint719_t(x : std_logic_vector) return uint719_t;
subtype int719_t is signed(718 downto 0);
constant int719_t_SLV_LEN : integer := 719;
function int719_t_to_slv(x : int719_t) return std_logic_vector;
function slv_to_int719_t(x : std_logic_vector) return int719_t;
subtype uint720_t is unsigned(719 downto 0);
constant uint720_t_SLV_LEN : integer := 720;
function uint720_t_to_slv(x : uint720_t) return std_logic_vector;
function slv_to_uint720_t(x : std_logic_vector) return uint720_t;
subtype int720_t is signed(719 downto 0);
constant int720_t_SLV_LEN : integer := 720;
function int720_t_to_slv(x : int720_t) return std_logic_vector;
function slv_to_int720_t(x : std_logic_vector) return int720_t;
subtype uint721_t is unsigned(720 downto 0);
constant uint721_t_SLV_LEN : integer := 721;
function uint721_t_to_slv(x : uint721_t) return std_logic_vector;
function slv_to_uint721_t(x : std_logic_vector) return uint721_t;
subtype int721_t is signed(720 downto 0);
constant int721_t_SLV_LEN : integer := 721;
function int721_t_to_slv(x : int721_t) return std_logic_vector;
function slv_to_int721_t(x : std_logic_vector) return int721_t;
subtype uint722_t is unsigned(721 downto 0);
constant uint722_t_SLV_LEN : integer := 722;
function uint722_t_to_slv(x : uint722_t) return std_logic_vector;
function slv_to_uint722_t(x : std_logic_vector) return uint722_t;
subtype int722_t is signed(721 downto 0);
constant int722_t_SLV_LEN : integer := 722;
function int722_t_to_slv(x : int722_t) return std_logic_vector;
function slv_to_int722_t(x : std_logic_vector) return int722_t;
subtype uint723_t is unsigned(722 downto 0);
constant uint723_t_SLV_LEN : integer := 723;
function uint723_t_to_slv(x : uint723_t) return std_logic_vector;
function slv_to_uint723_t(x : std_logic_vector) return uint723_t;
subtype int723_t is signed(722 downto 0);
constant int723_t_SLV_LEN : integer := 723;
function int723_t_to_slv(x : int723_t) return std_logic_vector;
function slv_to_int723_t(x : std_logic_vector) return int723_t;
subtype uint724_t is unsigned(723 downto 0);
constant uint724_t_SLV_LEN : integer := 724;
function uint724_t_to_slv(x : uint724_t) return std_logic_vector;
function slv_to_uint724_t(x : std_logic_vector) return uint724_t;
subtype int724_t is signed(723 downto 0);
constant int724_t_SLV_LEN : integer := 724;
function int724_t_to_slv(x : int724_t) return std_logic_vector;
function slv_to_int724_t(x : std_logic_vector) return int724_t;
subtype uint725_t is unsigned(724 downto 0);
constant uint725_t_SLV_LEN : integer := 725;
function uint725_t_to_slv(x : uint725_t) return std_logic_vector;
function slv_to_uint725_t(x : std_logic_vector) return uint725_t;
subtype int725_t is signed(724 downto 0);
constant int725_t_SLV_LEN : integer := 725;
function int725_t_to_slv(x : int725_t) return std_logic_vector;
function slv_to_int725_t(x : std_logic_vector) return int725_t;
subtype uint726_t is unsigned(725 downto 0);
constant uint726_t_SLV_LEN : integer := 726;
function uint726_t_to_slv(x : uint726_t) return std_logic_vector;
function slv_to_uint726_t(x : std_logic_vector) return uint726_t;
subtype int726_t is signed(725 downto 0);
constant int726_t_SLV_LEN : integer := 726;
function int726_t_to_slv(x : int726_t) return std_logic_vector;
function slv_to_int726_t(x : std_logic_vector) return int726_t;
subtype uint727_t is unsigned(726 downto 0);
constant uint727_t_SLV_LEN : integer := 727;
function uint727_t_to_slv(x : uint727_t) return std_logic_vector;
function slv_to_uint727_t(x : std_logic_vector) return uint727_t;
subtype int727_t is signed(726 downto 0);
constant int727_t_SLV_LEN : integer := 727;
function int727_t_to_slv(x : int727_t) return std_logic_vector;
function slv_to_int727_t(x : std_logic_vector) return int727_t;
subtype uint728_t is unsigned(727 downto 0);
constant uint728_t_SLV_LEN : integer := 728;
function uint728_t_to_slv(x : uint728_t) return std_logic_vector;
function slv_to_uint728_t(x : std_logic_vector) return uint728_t;
subtype int728_t is signed(727 downto 0);
constant int728_t_SLV_LEN : integer := 728;
function int728_t_to_slv(x : int728_t) return std_logic_vector;
function slv_to_int728_t(x : std_logic_vector) return int728_t;
subtype uint729_t is unsigned(728 downto 0);
constant uint729_t_SLV_LEN : integer := 729;
function uint729_t_to_slv(x : uint729_t) return std_logic_vector;
function slv_to_uint729_t(x : std_logic_vector) return uint729_t;
subtype int729_t is signed(728 downto 0);
constant int729_t_SLV_LEN : integer := 729;
function int729_t_to_slv(x : int729_t) return std_logic_vector;
function slv_to_int729_t(x : std_logic_vector) return int729_t;
subtype uint730_t is unsigned(729 downto 0);
constant uint730_t_SLV_LEN : integer := 730;
function uint730_t_to_slv(x : uint730_t) return std_logic_vector;
function slv_to_uint730_t(x : std_logic_vector) return uint730_t;
subtype int730_t is signed(729 downto 0);
constant int730_t_SLV_LEN : integer := 730;
function int730_t_to_slv(x : int730_t) return std_logic_vector;
function slv_to_int730_t(x : std_logic_vector) return int730_t;
subtype uint731_t is unsigned(730 downto 0);
constant uint731_t_SLV_LEN : integer := 731;
function uint731_t_to_slv(x : uint731_t) return std_logic_vector;
function slv_to_uint731_t(x : std_logic_vector) return uint731_t;
subtype int731_t is signed(730 downto 0);
constant int731_t_SLV_LEN : integer := 731;
function int731_t_to_slv(x : int731_t) return std_logic_vector;
function slv_to_int731_t(x : std_logic_vector) return int731_t;
subtype uint732_t is unsigned(731 downto 0);
constant uint732_t_SLV_LEN : integer := 732;
function uint732_t_to_slv(x : uint732_t) return std_logic_vector;
function slv_to_uint732_t(x : std_logic_vector) return uint732_t;
subtype int732_t is signed(731 downto 0);
constant int732_t_SLV_LEN : integer := 732;
function int732_t_to_slv(x : int732_t) return std_logic_vector;
function slv_to_int732_t(x : std_logic_vector) return int732_t;
subtype uint733_t is unsigned(732 downto 0);
constant uint733_t_SLV_LEN : integer := 733;
function uint733_t_to_slv(x : uint733_t) return std_logic_vector;
function slv_to_uint733_t(x : std_logic_vector) return uint733_t;
subtype int733_t is signed(732 downto 0);
constant int733_t_SLV_LEN : integer := 733;
function int733_t_to_slv(x : int733_t) return std_logic_vector;
function slv_to_int733_t(x : std_logic_vector) return int733_t;
subtype uint734_t is unsigned(733 downto 0);
constant uint734_t_SLV_LEN : integer := 734;
function uint734_t_to_slv(x : uint734_t) return std_logic_vector;
function slv_to_uint734_t(x : std_logic_vector) return uint734_t;
subtype int734_t is signed(733 downto 0);
constant int734_t_SLV_LEN : integer := 734;
function int734_t_to_slv(x : int734_t) return std_logic_vector;
function slv_to_int734_t(x : std_logic_vector) return int734_t;
subtype uint735_t is unsigned(734 downto 0);
constant uint735_t_SLV_LEN : integer := 735;
function uint735_t_to_slv(x : uint735_t) return std_logic_vector;
function slv_to_uint735_t(x : std_logic_vector) return uint735_t;
subtype int735_t is signed(734 downto 0);
constant int735_t_SLV_LEN : integer := 735;
function int735_t_to_slv(x : int735_t) return std_logic_vector;
function slv_to_int735_t(x : std_logic_vector) return int735_t;
subtype uint736_t is unsigned(735 downto 0);
constant uint736_t_SLV_LEN : integer := 736;
function uint736_t_to_slv(x : uint736_t) return std_logic_vector;
function slv_to_uint736_t(x : std_logic_vector) return uint736_t;
subtype int736_t is signed(735 downto 0);
constant int736_t_SLV_LEN : integer := 736;
function int736_t_to_slv(x : int736_t) return std_logic_vector;
function slv_to_int736_t(x : std_logic_vector) return int736_t;
subtype uint737_t is unsigned(736 downto 0);
constant uint737_t_SLV_LEN : integer := 737;
function uint737_t_to_slv(x : uint737_t) return std_logic_vector;
function slv_to_uint737_t(x : std_logic_vector) return uint737_t;
subtype int737_t is signed(736 downto 0);
constant int737_t_SLV_LEN : integer := 737;
function int737_t_to_slv(x : int737_t) return std_logic_vector;
function slv_to_int737_t(x : std_logic_vector) return int737_t;
subtype uint738_t is unsigned(737 downto 0);
constant uint738_t_SLV_LEN : integer := 738;
function uint738_t_to_slv(x : uint738_t) return std_logic_vector;
function slv_to_uint738_t(x : std_logic_vector) return uint738_t;
subtype int738_t is signed(737 downto 0);
constant int738_t_SLV_LEN : integer := 738;
function int738_t_to_slv(x : int738_t) return std_logic_vector;
function slv_to_int738_t(x : std_logic_vector) return int738_t;
subtype uint739_t is unsigned(738 downto 0);
constant uint739_t_SLV_LEN : integer := 739;
function uint739_t_to_slv(x : uint739_t) return std_logic_vector;
function slv_to_uint739_t(x : std_logic_vector) return uint739_t;
subtype int739_t is signed(738 downto 0);
constant int739_t_SLV_LEN : integer := 739;
function int739_t_to_slv(x : int739_t) return std_logic_vector;
function slv_to_int739_t(x : std_logic_vector) return int739_t;
subtype uint740_t is unsigned(739 downto 0);
constant uint740_t_SLV_LEN : integer := 740;
function uint740_t_to_slv(x : uint740_t) return std_logic_vector;
function slv_to_uint740_t(x : std_logic_vector) return uint740_t;
subtype int740_t is signed(739 downto 0);
constant int740_t_SLV_LEN : integer := 740;
function int740_t_to_slv(x : int740_t) return std_logic_vector;
function slv_to_int740_t(x : std_logic_vector) return int740_t;
subtype uint741_t is unsigned(740 downto 0);
constant uint741_t_SLV_LEN : integer := 741;
function uint741_t_to_slv(x : uint741_t) return std_logic_vector;
function slv_to_uint741_t(x : std_logic_vector) return uint741_t;
subtype int741_t is signed(740 downto 0);
constant int741_t_SLV_LEN : integer := 741;
function int741_t_to_slv(x : int741_t) return std_logic_vector;
function slv_to_int741_t(x : std_logic_vector) return int741_t;
subtype uint742_t is unsigned(741 downto 0);
constant uint742_t_SLV_LEN : integer := 742;
function uint742_t_to_slv(x : uint742_t) return std_logic_vector;
function slv_to_uint742_t(x : std_logic_vector) return uint742_t;
subtype int742_t is signed(741 downto 0);
constant int742_t_SLV_LEN : integer := 742;
function int742_t_to_slv(x : int742_t) return std_logic_vector;
function slv_to_int742_t(x : std_logic_vector) return int742_t;
subtype uint743_t is unsigned(742 downto 0);
constant uint743_t_SLV_LEN : integer := 743;
function uint743_t_to_slv(x : uint743_t) return std_logic_vector;
function slv_to_uint743_t(x : std_logic_vector) return uint743_t;
subtype int743_t is signed(742 downto 0);
constant int743_t_SLV_LEN : integer := 743;
function int743_t_to_slv(x : int743_t) return std_logic_vector;
function slv_to_int743_t(x : std_logic_vector) return int743_t;
subtype uint744_t is unsigned(743 downto 0);
constant uint744_t_SLV_LEN : integer := 744;
function uint744_t_to_slv(x : uint744_t) return std_logic_vector;
function slv_to_uint744_t(x : std_logic_vector) return uint744_t;
subtype int744_t is signed(743 downto 0);
constant int744_t_SLV_LEN : integer := 744;
function int744_t_to_slv(x : int744_t) return std_logic_vector;
function slv_to_int744_t(x : std_logic_vector) return int744_t;
subtype uint745_t is unsigned(744 downto 0);
constant uint745_t_SLV_LEN : integer := 745;
function uint745_t_to_slv(x : uint745_t) return std_logic_vector;
function slv_to_uint745_t(x : std_logic_vector) return uint745_t;
subtype int745_t is signed(744 downto 0);
constant int745_t_SLV_LEN : integer := 745;
function int745_t_to_slv(x : int745_t) return std_logic_vector;
function slv_to_int745_t(x : std_logic_vector) return int745_t;
subtype uint746_t is unsigned(745 downto 0);
constant uint746_t_SLV_LEN : integer := 746;
function uint746_t_to_slv(x : uint746_t) return std_logic_vector;
function slv_to_uint746_t(x : std_logic_vector) return uint746_t;
subtype int746_t is signed(745 downto 0);
constant int746_t_SLV_LEN : integer := 746;
function int746_t_to_slv(x : int746_t) return std_logic_vector;
function slv_to_int746_t(x : std_logic_vector) return int746_t;
subtype uint747_t is unsigned(746 downto 0);
constant uint747_t_SLV_LEN : integer := 747;
function uint747_t_to_slv(x : uint747_t) return std_logic_vector;
function slv_to_uint747_t(x : std_logic_vector) return uint747_t;
subtype int747_t is signed(746 downto 0);
constant int747_t_SLV_LEN : integer := 747;
function int747_t_to_slv(x : int747_t) return std_logic_vector;
function slv_to_int747_t(x : std_logic_vector) return int747_t;
subtype uint748_t is unsigned(747 downto 0);
constant uint748_t_SLV_LEN : integer := 748;
function uint748_t_to_slv(x : uint748_t) return std_logic_vector;
function slv_to_uint748_t(x : std_logic_vector) return uint748_t;
subtype int748_t is signed(747 downto 0);
constant int748_t_SLV_LEN : integer := 748;
function int748_t_to_slv(x : int748_t) return std_logic_vector;
function slv_to_int748_t(x : std_logic_vector) return int748_t;
subtype uint749_t is unsigned(748 downto 0);
constant uint749_t_SLV_LEN : integer := 749;
function uint749_t_to_slv(x : uint749_t) return std_logic_vector;
function slv_to_uint749_t(x : std_logic_vector) return uint749_t;
subtype int749_t is signed(748 downto 0);
constant int749_t_SLV_LEN : integer := 749;
function int749_t_to_slv(x : int749_t) return std_logic_vector;
function slv_to_int749_t(x : std_logic_vector) return int749_t;
subtype uint750_t is unsigned(749 downto 0);
constant uint750_t_SLV_LEN : integer := 750;
function uint750_t_to_slv(x : uint750_t) return std_logic_vector;
function slv_to_uint750_t(x : std_logic_vector) return uint750_t;
subtype int750_t is signed(749 downto 0);
constant int750_t_SLV_LEN : integer := 750;
function int750_t_to_slv(x : int750_t) return std_logic_vector;
function slv_to_int750_t(x : std_logic_vector) return int750_t;
subtype uint751_t is unsigned(750 downto 0);
constant uint751_t_SLV_LEN : integer := 751;
function uint751_t_to_slv(x : uint751_t) return std_logic_vector;
function slv_to_uint751_t(x : std_logic_vector) return uint751_t;
subtype int751_t is signed(750 downto 0);
constant int751_t_SLV_LEN : integer := 751;
function int751_t_to_slv(x : int751_t) return std_logic_vector;
function slv_to_int751_t(x : std_logic_vector) return int751_t;
subtype uint752_t is unsigned(751 downto 0);
constant uint752_t_SLV_LEN : integer := 752;
function uint752_t_to_slv(x : uint752_t) return std_logic_vector;
function slv_to_uint752_t(x : std_logic_vector) return uint752_t;
subtype int752_t is signed(751 downto 0);
constant int752_t_SLV_LEN : integer := 752;
function int752_t_to_slv(x : int752_t) return std_logic_vector;
function slv_to_int752_t(x : std_logic_vector) return int752_t;
subtype uint753_t is unsigned(752 downto 0);
constant uint753_t_SLV_LEN : integer := 753;
function uint753_t_to_slv(x : uint753_t) return std_logic_vector;
function slv_to_uint753_t(x : std_logic_vector) return uint753_t;
subtype int753_t is signed(752 downto 0);
constant int753_t_SLV_LEN : integer := 753;
function int753_t_to_slv(x : int753_t) return std_logic_vector;
function slv_to_int753_t(x : std_logic_vector) return int753_t;
subtype uint754_t is unsigned(753 downto 0);
constant uint754_t_SLV_LEN : integer := 754;
function uint754_t_to_slv(x : uint754_t) return std_logic_vector;
function slv_to_uint754_t(x : std_logic_vector) return uint754_t;
subtype int754_t is signed(753 downto 0);
constant int754_t_SLV_LEN : integer := 754;
function int754_t_to_slv(x : int754_t) return std_logic_vector;
function slv_to_int754_t(x : std_logic_vector) return int754_t;
subtype uint755_t is unsigned(754 downto 0);
constant uint755_t_SLV_LEN : integer := 755;
function uint755_t_to_slv(x : uint755_t) return std_logic_vector;
function slv_to_uint755_t(x : std_logic_vector) return uint755_t;
subtype int755_t is signed(754 downto 0);
constant int755_t_SLV_LEN : integer := 755;
function int755_t_to_slv(x : int755_t) return std_logic_vector;
function slv_to_int755_t(x : std_logic_vector) return int755_t;
subtype uint756_t is unsigned(755 downto 0);
constant uint756_t_SLV_LEN : integer := 756;
function uint756_t_to_slv(x : uint756_t) return std_logic_vector;
function slv_to_uint756_t(x : std_logic_vector) return uint756_t;
subtype int756_t is signed(755 downto 0);
constant int756_t_SLV_LEN : integer := 756;
function int756_t_to_slv(x : int756_t) return std_logic_vector;
function slv_to_int756_t(x : std_logic_vector) return int756_t;
subtype uint757_t is unsigned(756 downto 0);
constant uint757_t_SLV_LEN : integer := 757;
function uint757_t_to_slv(x : uint757_t) return std_logic_vector;
function slv_to_uint757_t(x : std_logic_vector) return uint757_t;
subtype int757_t is signed(756 downto 0);
constant int757_t_SLV_LEN : integer := 757;
function int757_t_to_slv(x : int757_t) return std_logic_vector;
function slv_to_int757_t(x : std_logic_vector) return int757_t;
subtype uint758_t is unsigned(757 downto 0);
constant uint758_t_SLV_LEN : integer := 758;
function uint758_t_to_slv(x : uint758_t) return std_logic_vector;
function slv_to_uint758_t(x : std_logic_vector) return uint758_t;
subtype int758_t is signed(757 downto 0);
constant int758_t_SLV_LEN : integer := 758;
function int758_t_to_slv(x : int758_t) return std_logic_vector;
function slv_to_int758_t(x : std_logic_vector) return int758_t;
subtype uint759_t is unsigned(758 downto 0);
constant uint759_t_SLV_LEN : integer := 759;
function uint759_t_to_slv(x : uint759_t) return std_logic_vector;
function slv_to_uint759_t(x : std_logic_vector) return uint759_t;
subtype int759_t is signed(758 downto 0);
constant int759_t_SLV_LEN : integer := 759;
function int759_t_to_slv(x : int759_t) return std_logic_vector;
function slv_to_int759_t(x : std_logic_vector) return int759_t;
subtype uint760_t is unsigned(759 downto 0);
constant uint760_t_SLV_LEN : integer := 760;
function uint760_t_to_slv(x : uint760_t) return std_logic_vector;
function slv_to_uint760_t(x : std_logic_vector) return uint760_t;
subtype int760_t is signed(759 downto 0);
constant int760_t_SLV_LEN : integer := 760;
function int760_t_to_slv(x : int760_t) return std_logic_vector;
function slv_to_int760_t(x : std_logic_vector) return int760_t;
subtype uint761_t is unsigned(760 downto 0);
constant uint761_t_SLV_LEN : integer := 761;
function uint761_t_to_slv(x : uint761_t) return std_logic_vector;
function slv_to_uint761_t(x : std_logic_vector) return uint761_t;
subtype int761_t is signed(760 downto 0);
constant int761_t_SLV_LEN : integer := 761;
function int761_t_to_slv(x : int761_t) return std_logic_vector;
function slv_to_int761_t(x : std_logic_vector) return int761_t;
subtype uint762_t is unsigned(761 downto 0);
constant uint762_t_SLV_LEN : integer := 762;
function uint762_t_to_slv(x : uint762_t) return std_logic_vector;
function slv_to_uint762_t(x : std_logic_vector) return uint762_t;
subtype int762_t is signed(761 downto 0);
constant int762_t_SLV_LEN : integer := 762;
function int762_t_to_slv(x : int762_t) return std_logic_vector;
function slv_to_int762_t(x : std_logic_vector) return int762_t;
subtype uint763_t is unsigned(762 downto 0);
constant uint763_t_SLV_LEN : integer := 763;
function uint763_t_to_slv(x : uint763_t) return std_logic_vector;
function slv_to_uint763_t(x : std_logic_vector) return uint763_t;
subtype int763_t is signed(762 downto 0);
constant int763_t_SLV_LEN : integer := 763;
function int763_t_to_slv(x : int763_t) return std_logic_vector;
function slv_to_int763_t(x : std_logic_vector) return int763_t;
subtype uint764_t is unsigned(763 downto 0);
constant uint764_t_SLV_LEN : integer := 764;
function uint764_t_to_slv(x : uint764_t) return std_logic_vector;
function slv_to_uint764_t(x : std_logic_vector) return uint764_t;
subtype int764_t is signed(763 downto 0);
constant int764_t_SLV_LEN : integer := 764;
function int764_t_to_slv(x : int764_t) return std_logic_vector;
function slv_to_int764_t(x : std_logic_vector) return int764_t;
subtype uint765_t is unsigned(764 downto 0);
constant uint765_t_SLV_LEN : integer := 765;
function uint765_t_to_slv(x : uint765_t) return std_logic_vector;
function slv_to_uint765_t(x : std_logic_vector) return uint765_t;
subtype int765_t is signed(764 downto 0);
constant int765_t_SLV_LEN : integer := 765;
function int765_t_to_slv(x : int765_t) return std_logic_vector;
function slv_to_int765_t(x : std_logic_vector) return int765_t;
subtype uint766_t is unsigned(765 downto 0);
constant uint766_t_SLV_LEN : integer := 766;
function uint766_t_to_slv(x : uint766_t) return std_logic_vector;
function slv_to_uint766_t(x : std_logic_vector) return uint766_t;
subtype int766_t is signed(765 downto 0);
constant int766_t_SLV_LEN : integer := 766;
function int766_t_to_slv(x : int766_t) return std_logic_vector;
function slv_to_int766_t(x : std_logic_vector) return int766_t;
subtype uint767_t is unsigned(766 downto 0);
constant uint767_t_SLV_LEN : integer := 767;
function uint767_t_to_slv(x : uint767_t) return std_logic_vector;
function slv_to_uint767_t(x : std_logic_vector) return uint767_t;
subtype int767_t is signed(766 downto 0);
constant int767_t_SLV_LEN : integer := 767;
function int767_t_to_slv(x : int767_t) return std_logic_vector;
function slv_to_int767_t(x : std_logic_vector) return int767_t;
subtype uint768_t is unsigned(767 downto 0);
constant uint768_t_SLV_LEN : integer := 768;
function uint768_t_to_slv(x : uint768_t) return std_logic_vector;
function slv_to_uint768_t(x : std_logic_vector) return uint768_t;
subtype int768_t is signed(767 downto 0);
constant int768_t_SLV_LEN : integer := 768;
function int768_t_to_slv(x : int768_t) return std_logic_vector;
function slv_to_int768_t(x : std_logic_vector) return int768_t;
subtype uint769_t is unsigned(768 downto 0);
constant uint769_t_SLV_LEN : integer := 769;
function uint769_t_to_slv(x : uint769_t) return std_logic_vector;
function slv_to_uint769_t(x : std_logic_vector) return uint769_t;
subtype int769_t is signed(768 downto 0);
constant int769_t_SLV_LEN : integer := 769;
function int769_t_to_slv(x : int769_t) return std_logic_vector;
function slv_to_int769_t(x : std_logic_vector) return int769_t;
subtype uint770_t is unsigned(769 downto 0);
constant uint770_t_SLV_LEN : integer := 770;
function uint770_t_to_slv(x : uint770_t) return std_logic_vector;
function slv_to_uint770_t(x : std_logic_vector) return uint770_t;
subtype int770_t is signed(769 downto 0);
constant int770_t_SLV_LEN : integer := 770;
function int770_t_to_slv(x : int770_t) return std_logic_vector;
function slv_to_int770_t(x : std_logic_vector) return int770_t;
subtype uint771_t is unsigned(770 downto 0);
constant uint771_t_SLV_LEN : integer := 771;
function uint771_t_to_slv(x : uint771_t) return std_logic_vector;
function slv_to_uint771_t(x : std_logic_vector) return uint771_t;
subtype int771_t is signed(770 downto 0);
constant int771_t_SLV_LEN : integer := 771;
function int771_t_to_slv(x : int771_t) return std_logic_vector;
function slv_to_int771_t(x : std_logic_vector) return int771_t;
subtype uint772_t is unsigned(771 downto 0);
constant uint772_t_SLV_LEN : integer := 772;
function uint772_t_to_slv(x : uint772_t) return std_logic_vector;
function slv_to_uint772_t(x : std_logic_vector) return uint772_t;
subtype int772_t is signed(771 downto 0);
constant int772_t_SLV_LEN : integer := 772;
function int772_t_to_slv(x : int772_t) return std_logic_vector;
function slv_to_int772_t(x : std_logic_vector) return int772_t;
subtype uint773_t is unsigned(772 downto 0);
constant uint773_t_SLV_LEN : integer := 773;
function uint773_t_to_slv(x : uint773_t) return std_logic_vector;
function slv_to_uint773_t(x : std_logic_vector) return uint773_t;
subtype int773_t is signed(772 downto 0);
constant int773_t_SLV_LEN : integer := 773;
function int773_t_to_slv(x : int773_t) return std_logic_vector;
function slv_to_int773_t(x : std_logic_vector) return int773_t;
subtype uint774_t is unsigned(773 downto 0);
constant uint774_t_SLV_LEN : integer := 774;
function uint774_t_to_slv(x : uint774_t) return std_logic_vector;
function slv_to_uint774_t(x : std_logic_vector) return uint774_t;
subtype int774_t is signed(773 downto 0);
constant int774_t_SLV_LEN : integer := 774;
function int774_t_to_slv(x : int774_t) return std_logic_vector;
function slv_to_int774_t(x : std_logic_vector) return int774_t;
subtype uint775_t is unsigned(774 downto 0);
constant uint775_t_SLV_LEN : integer := 775;
function uint775_t_to_slv(x : uint775_t) return std_logic_vector;
function slv_to_uint775_t(x : std_logic_vector) return uint775_t;
subtype int775_t is signed(774 downto 0);
constant int775_t_SLV_LEN : integer := 775;
function int775_t_to_slv(x : int775_t) return std_logic_vector;
function slv_to_int775_t(x : std_logic_vector) return int775_t;
subtype uint776_t is unsigned(775 downto 0);
constant uint776_t_SLV_LEN : integer := 776;
function uint776_t_to_slv(x : uint776_t) return std_logic_vector;
function slv_to_uint776_t(x : std_logic_vector) return uint776_t;
subtype int776_t is signed(775 downto 0);
constant int776_t_SLV_LEN : integer := 776;
function int776_t_to_slv(x : int776_t) return std_logic_vector;
function slv_to_int776_t(x : std_logic_vector) return int776_t;
subtype uint777_t is unsigned(776 downto 0);
constant uint777_t_SLV_LEN : integer := 777;
function uint777_t_to_slv(x : uint777_t) return std_logic_vector;
function slv_to_uint777_t(x : std_logic_vector) return uint777_t;
subtype int777_t is signed(776 downto 0);
constant int777_t_SLV_LEN : integer := 777;
function int777_t_to_slv(x : int777_t) return std_logic_vector;
function slv_to_int777_t(x : std_logic_vector) return int777_t;
subtype uint778_t is unsigned(777 downto 0);
constant uint778_t_SLV_LEN : integer := 778;
function uint778_t_to_slv(x : uint778_t) return std_logic_vector;
function slv_to_uint778_t(x : std_logic_vector) return uint778_t;
subtype int778_t is signed(777 downto 0);
constant int778_t_SLV_LEN : integer := 778;
function int778_t_to_slv(x : int778_t) return std_logic_vector;
function slv_to_int778_t(x : std_logic_vector) return int778_t;
subtype uint779_t is unsigned(778 downto 0);
constant uint779_t_SLV_LEN : integer := 779;
function uint779_t_to_slv(x : uint779_t) return std_logic_vector;
function slv_to_uint779_t(x : std_logic_vector) return uint779_t;
subtype int779_t is signed(778 downto 0);
constant int779_t_SLV_LEN : integer := 779;
function int779_t_to_slv(x : int779_t) return std_logic_vector;
function slv_to_int779_t(x : std_logic_vector) return int779_t;
subtype uint780_t is unsigned(779 downto 0);
constant uint780_t_SLV_LEN : integer := 780;
function uint780_t_to_slv(x : uint780_t) return std_logic_vector;
function slv_to_uint780_t(x : std_logic_vector) return uint780_t;
subtype int780_t is signed(779 downto 0);
constant int780_t_SLV_LEN : integer := 780;
function int780_t_to_slv(x : int780_t) return std_logic_vector;
function slv_to_int780_t(x : std_logic_vector) return int780_t;
subtype uint781_t is unsigned(780 downto 0);
constant uint781_t_SLV_LEN : integer := 781;
function uint781_t_to_slv(x : uint781_t) return std_logic_vector;
function slv_to_uint781_t(x : std_logic_vector) return uint781_t;
subtype int781_t is signed(780 downto 0);
constant int781_t_SLV_LEN : integer := 781;
function int781_t_to_slv(x : int781_t) return std_logic_vector;
function slv_to_int781_t(x : std_logic_vector) return int781_t;
subtype uint782_t is unsigned(781 downto 0);
constant uint782_t_SLV_LEN : integer := 782;
function uint782_t_to_slv(x : uint782_t) return std_logic_vector;
function slv_to_uint782_t(x : std_logic_vector) return uint782_t;
subtype int782_t is signed(781 downto 0);
constant int782_t_SLV_LEN : integer := 782;
function int782_t_to_slv(x : int782_t) return std_logic_vector;
function slv_to_int782_t(x : std_logic_vector) return int782_t;
subtype uint783_t is unsigned(782 downto 0);
constant uint783_t_SLV_LEN : integer := 783;
function uint783_t_to_slv(x : uint783_t) return std_logic_vector;
function slv_to_uint783_t(x : std_logic_vector) return uint783_t;
subtype int783_t is signed(782 downto 0);
constant int783_t_SLV_LEN : integer := 783;
function int783_t_to_slv(x : int783_t) return std_logic_vector;
function slv_to_int783_t(x : std_logic_vector) return int783_t;
subtype uint784_t is unsigned(783 downto 0);
constant uint784_t_SLV_LEN : integer := 784;
function uint784_t_to_slv(x : uint784_t) return std_logic_vector;
function slv_to_uint784_t(x : std_logic_vector) return uint784_t;
subtype int784_t is signed(783 downto 0);
constant int784_t_SLV_LEN : integer := 784;
function int784_t_to_slv(x : int784_t) return std_logic_vector;
function slv_to_int784_t(x : std_logic_vector) return int784_t;
subtype uint785_t is unsigned(784 downto 0);
constant uint785_t_SLV_LEN : integer := 785;
function uint785_t_to_slv(x : uint785_t) return std_logic_vector;
function slv_to_uint785_t(x : std_logic_vector) return uint785_t;
subtype int785_t is signed(784 downto 0);
constant int785_t_SLV_LEN : integer := 785;
function int785_t_to_slv(x : int785_t) return std_logic_vector;
function slv_to_int785_t(x : std_logic_vector) return int785_t;
subtype uint786_t is unsigned(785 downto 0);
constant uint786_t_SLV_LEN : integer := 786;
function uint786_t_to_slv(x : uint786_t) return std_logic_vector;
function slv_to_uint786_t(x : std_logic_vector) return uint786_t;
subtype int786_t is signed(785 downto 0);
constant int786_t_SLV_LEN : integer := 786;
function int786_t_to_slv(x : int786_t) return std_logic_vector;
function slv_to_int786_t(x : std_logic_vector) return int786_t;
subtype uint787_t is unsigned(786 downto 0);
constant uint787_t_SLV_LEN : integer := 787;
function uint787_t_to_slv(x : uint787_t) return std_logic_vector;
function slv_to_uint787_t(x : std_logic_vector) return uint787_t;
subtype int787_t is signed(786 downto 0);
constant int787_t_SLV_LEN : integer := 787;
function int787_t_to_slv(x : int787_t) return std_logic_vector;
function slv_to_int787_t(x : std_logic_vector) return int787_t;
subtype uint788_t is unsigned(787 downto 0);
constant uint788_t_SLV_LEN : integer := 788;
function uint788_t_to_slv(x : uint788_t) return std_logic_vector;
function slv_to_uint788_t(x : std_logic_vector) return uint788_t;
subtype int788_t is signed(787 downto 0);
constant int788_t_SLV_LEN : integer := 788;
function int788_t_to_slv(x : int788_t) return std_logic_vector;
function slv_to_int788_t(x : std_logic_vector) return int788_t;
subtype uint789_t is unsigned(788 downto 0);
constant uint789_t_SLV_LEN : integer := 789;
function uint789_t_to_slv(x : uint789_t) return std_logic_vector;
function slv_to_uint789_t(x : std_logic_vector) return uint789_t;
subtype int789_t is signed(788 downto 0);
constant int789_t_SLV_LEN : integer := 789;
function int789_t_to_slv(x : int789_t) return std_logic_vector;
function slv_to_int789_t(x : std_logic_vector) return int789_t;
subtype uint790_t is unsigned(789 downto 0);
constant uint790_t_SLV_LEN : integer := 790;
function uint790_t_to_slv(x : uint790_t) return std_logic_vector;
function slv_to_uint790_t(x : std_logic_vector) return uint790_t;
subtype int790_t is signed(789 downto 0);
constant int790_t_SLV_LEN : integer := 790;
function int790_t_to_slv(x : int790_t) return std_logic_vector;
function slv_to_int790_t(x : std_logic_vector) return int790_t;
subtype uint791_t is unsigned(790 downto 0);
constant uint791_t_SLV_LEN : integer := 791;
function uint791_t_to_slv(x : uint791_t) return std_logic_vector;
function slv_to_uint791_t(x : std_logic_vector) return uint791_t;
subtype int791_t is signed(790 downto 0);
constant int791_t_SLV_LEN : integer := 791;
function int791_t_to_slv(x : int791_t) return std_logic_vector;
function slv_to_int791_t(x : std_logic_vector) return int791_t;
subtype uint792_t is unsigned(791 downto 0);
constant uint792_t_SLV_LEN : integer := 792;
function uint792_t_to_slv(x : uint792_t) return std_logic_vector;
function slv_to_uint792_t(x : std_logic_vector) return uint792_t;
subtype int792_t is signed(791 downto 0);
constant int792_t_SLV_LEN : integer := 792;
function int792_t_to_slv(x : int792_t) return std_logic_vector;
function slv_to_int792_t(x : std_logic_vector) return int792_t;
subtype uint793_t is unsigned(792 downto 0);
constant uint793_t_SLV_LEN : integer := 793;
function uint793_t_to_slv(x : uint793_t) return std_logic_vector;
function slv_to_uint793_t(x : std_logic_vector) return uint793_t;
subtype int793_t is signed(792 downto 0);
constant int793_t_SLV_LEN : integer := 793;
function int793_t_to_slv(x : int793_t) return std_logic_vector;
function slv_to_int793_t(x : std_logic_vector) return int793_t;
subtype uint794_t is unsigned(793 downto 0);
constant uint794_t_SLV_LEN : integer := 794;
function uint794_t_to_slv(x : uint794_t) return std_logic_vector;
function slv_to_uint794_t(x : std_logic_vector) return uint794_t;
subtype int794_t is signed(793 downto 0);
constant int794_t_SLV_LEN : integer := 794;
function int794_t_to_slv(x : int794_t) return std_logic_vector;
function slv_to_int794_t(x : std_logic_vector) return int794_t;
subtype uint795_t is unsigned(794 downto 0);
constant uint795_t_SLV_LEN : integer := 795;
function uint795_t_to_slv(x : uint795_t) return std_logic_vector;
function slv_to_uint795_t(x : std_logic_vector) return uint795_t;
subtype int795_t is signed(794 downto 0);
constant int795_t_SLV_LEN : integer := 795;
function int795_t_to_slv(x : int795_t) return std_logic_vector;
function slv_to_int795_t(x : std_logic_vector) return int795_t;
subtype uint796_t is unsigned(795 downto 0);
constant uint796_t_SLV_LEN : integer := 796;
function uint796_t_to_slv(x : uint796_t) return std_logic_vector;
function slv_to_uint796_t(x : std_logic_vector) return uint796_t;
subtype int796_t is signed(795 downto 0);
constant int796_t_SLV_LEN : integer := 796;
function int796_t_to_slv(x : int796_t) return std_logic_vector;
function slv_to_int796_t(x : std_logic_vector) return int796_t;
subtype uint797_t is unsigned(796 downto 0);
constant uint797_t_SLV_LEN : integer := 797;
function uint797_t_to_slv(x : uint797_t) return std_logic_vector;
function slv_to_uint797_t(x : std_logic_vector) return uint797_t;
subtype int797_t is signed(796 downto 0);
constant int797_t_SLV_LEN : integer := 797;
function int797_t_to_slv(x : int797_t) return std_logic_vector;
function slv_to_int797_t(x : std_logic_vector) return int797_t;
subtype uint798_t is unsigned(797 downto 0);
constant uint798_t_SLV_LEN : integer := 798;
function uint798_t_to_slv(x : uint798_t) return std_logic_vector;
function slv_to_uint798_t(x : std_logic_vector) return uint798_t;
subtype int798_t is signed(797 downto 0);
constant int798_t_SLV_LEN : integer := 798;
function int798_t_to_slv(x : int798_t) return std_logic_vector;
function slv_to_int798_t(x : std_logic_vector) return int798_t;
subtype uint799_t is unsigned(798 downto 0);
constant uint799_t_SLV_LEN : integer := 799;
function uint799_t_to_slv(x : uint799_t) return std_logic_vector;
function slv_to_uint799_t(x : std_logic_vector) return uint799_t;
subtype int799_t is signed(798 downto 0);
constant int799_t_SLV_LEN : integer := 799;
function int799_t_to_slv(x : int799_t) return std_logic_vector;
function slv_to_int799_t(x : std_logic_vector) return int799_t;
subtype uint800_t is unsigned(799 downto 0);
constant uint800_t_SLV_LEN : integer := 800;
function uint800_t_to_slv(x : uint800_t) return std_logic_vector;
function slv_to_uint800_t(x : std_logic_vector) return uint800_t;
subtype int800_t is signed(799 downto 0);
constant int800_t_SLV_LEN : integer := 800;
function int800_t_to_slv(x : int800_t) return std_logic_vector;
function slv_to_int800_t(x : std_logic_vector) return int800_t;
subtype uint801_t is unsigned(800 downto 0);
constant uint801_t_SLV_LEN : integer := 801;
function uint801_t_to_slv(x : uint801_t) return std_logic_vector;
function slv_to_uint801_t(x : std_logic_vector) return uint801_t;
subtype int801_t is signed(800 downto 0);
constant int801_t_SLV_LEN : integer := 801;
function int801_t_to_slv(x : int801_t) return std_logic_vector;
function slv_to_int801_t(x : std_logic_vector) return int801_t;
subtype uint802_t is unsigned(801 downto 0);
constant uint802_t_SLV_LEN : integer := 802;
function uint802_t_to_slv(x : uint802_t) return std_logic_vector;
function slv_to_uint802_t(x : std_logic_vector) return uint802_t;
subtype int802_t is signed(801 downto 0);
constant int802_t_SLV_LEN : integer := 802;
function int802_t_to_slv(x : int802_t) return std_logic_vector;
function slv_to_int802_t(x : std_logic_vector) return int802_t;
subtype uint803_t is unsigned(802 downto 0);
constant uint803_t_SLV_LEN : integer := 803;
function uint803_t_to_slv(x : uint803_t) return std_logic_vector;
function slv_to_uint803_t(x : std_logic_vector) return uint803_t;
subtype int803_t is signed(802 downto 0);
constant int803_t_SLV_LEN : integer := 803;
function int803_t_to_slv(x : int803_t) return std_logic_vector;
function slv_to_int803_t(x : std_logic_vector) return int803_t;
subtype uint804_t is unsigned(803 downto 0);
constant uint804_t_SLV_LEN : integer := 804;
function uint804_t_to_slv(x : uint804_t) return std_logic_vector;
function slv_to_uint804_t(x : std_logic_vector) return uint804_t;
subtype int804_t is signed(803 downto 0);
constant int804_t_SLV_LEN : integer := 804;
function int804_t_to_slv(x : int804_t) return std_logic_vector;
function slv_to_int804_t(x : std_logic_vector) return int804_t;
subtype uint805_t is unsigned(804 downto 0);
constant uint805_t_SLV_LEN : integer := 805;
function uint805_t_to_slv(x : uint805_t) return std_logic_vector;
function slv_to_uint805_t(x : std_logic_vector) return uint805_t;
subtype int805_t is signed(804 downto 0);
constant int805_t_SLV_LEN : integer := 805;
function int805_t_to_slv(x : int805_t) return std_logic_vector;
function slv_to_int805_t(x : std_logic_vector) return int805_t;
subtype uint806_t is unsigned(805 downto 0);
constant uint806_t_SLV_LEN : integer := 806;
function uint806_t_to_slv(x : uint806_t) return std_logic_vector;
function slv_to_uint806_t(x : std_logic_vector) return uint806_t;
subtype int806_t is signed(805 downto 0);
constant int806_t_SLV_LEN : integer := 806;
function int806_t_to_slv(x : int806_t) return std_logic_vector;
function slv_to_int806_t(x : std_logic_vector) return int806_t;
subtype uint807_t is unsigned(806 downto 0);
constant uint807_t_SLV_LEN : integer := 807;
function uint807_t_to_slv(x : uint807_t) return std_logic_vector;
function slv_to_uint807_t(x : std_logic_vector) return uint807_t;
subtype int807_t is signed(806 downto 0);
constant int807_t_SLV_LEN : integer := 807;
function int807_t_to_slv(x : int807_t) return std_logic_vector;
function slv_to_int807_t(x : std_logic_vector) return int807_t;
subtype uint808_t is unsigned(807 downto 0);
constant uint808_t_SLV_LEN : integer := 808;
function uint808_t_to_slv(x : uint808_t) return std_logic_vector;
function slv_to_uint808_t(x : std_logic_vector) return uint808_t;
subtype int808_t is signed(807 downto 0);
constant int808_t_SLV_LEN : integer := 808;
function int808_t_to_slv(x : int808_t) return std_logic_vector;
function slv_to_int808_t(x : std_logic_vector) return int808_t;
subtype uint809_t is unsigned(808 downto 0);
constant uint809_t_SLV_LEN : integer := 809;
function uint809_t_to_slv(x : uint809_t) return std_logic_vector;
function slv_to_uint809_t(x : std_logic_vector) return uint809_t;
subtype int809_t is signed(808 downto 0);
constant int809_t_SLV_LEN : integer := 809;
function int809_t_to_slv(x : int809_t) return std_logic_vector;
function slv_to_int809_t(x : std_logic_vector) return int809_t;
subtype uint810_t is unsigned(809 downto 0);
constant uint810_t_SLV_LEN : integer := 810;
function uint810_t_to_slv(x : uint810_t) return std_logic_vector;
function slv_to_uint810_t(x : std_logic_vector) return uint810_t;
subtype int810_t is signed(809 downto 0);
constant int810_t_SLV_LEN : integer := 810;
function int810_t_to_slv(x : int810_t) return std_logic_vector;
function slv_to_int810_t(x : std_logic_vector) return int810_t;
subtype uint811_t is unsigned(810 downto 0);
constant uint811_t_SLV_LEN : integer := 811;
function uint811_t_to_slv(x : uint811_t) return std_logic_vector;
function slv_to_uint811_t(x : std_logic_vector) return uint811_t;
subtype int811_t is signed(810 downto 0);
constant int811_t_SLV_LEN : integer := 811;
function int811_t_to_slv(x : int811_t) return std_logic_vector;
function slv_to_int811_t(x : std_logic_vector) return int811_t;
subtype uint812_t is unsigned(811 downto 0);
constant uint812_t_SLV_LEN : integer := 812;
function uint812_t_to_slv(x : uint812_t) return std_logic_vector;
function slv_to_uint812_t(x : std_logic_vector) return uint812_t;
subtype int812_t is signed(811 downto 0);
constant int812_t_SLV_LEN : integer := 812;
function int812_t_to_slv(x : int812_t) return std_logic_vector;
function slv_to_int812_t(x : std_logic_vector) return int812_t;
subtype uint813_t is unsigned(812 downto 0);
constant uint813_t_SLV_LEN : integer := 813;
function uint813_t_to_slv(x : uint813_t) return std_logic_vector;
function slv_to_uint813_t(x : std_logic_vector) return uint813_t;
subtype int813_t is signed(812 downto 0);
constant int813_t_SLV_LEN : integer := 813;
function int813_t_to_slv(x : int813_t) return std_logic_vector;
function slv_to_int813_t(x : std_logic_vector) return int813_t;
subtype uint814_t is unsigned(813 downto 0);
constant uint814_t_SLV_LEN : integer := 814;
function uint814_t_to_slv(x : uint814_t) return std_logic_vector;
function slv_to_uint814_t(x : std_logic_vector) return uint814_t;
subtype int814_t is signed(813 downto 0);
constant int814_t_SLV_LEN : integer := 814;
function int814_t_to_slv(x : int814_t) return std_logic_vector;
function slv_to_int814_t(x : std_logic_vector) return int814_t;
subtype uint815_t is unsigned(814 downto 0);
constant uint815_t_SLV_LEN : integer := 815;
function uint815_t_to_slv(x : uint815_t) return std_logic_vector;
function slv_to_uint815_t(x : std_logic_vector) return uint815_t;
subtype int815_t is signed(814 downto 0);
constant int815_t_SLV_LEN : integer := 815;
function int815_t_to_slv(x : int815_t) return std_logic_vector;
function slv_to_int815_t(x : std_logic_vector) return int815_t;
subtype uint816_t is unsigned(815 downto 0);
constant uint816_t_SLV_LEN : integer := 816;
function uint816_t_to_slv(x : uint816_t) return std_logic_vector;
function slv_to_uint816_t(x : std_logic_vector) return uint816_t;
subtype int816_t is signed(815 downto 0);
constant int816_t_SLV_LEN : integer := 816;
function int816_t_to_slv(x : int816_t) return std_logic_vector;
function slv_to_int816_t(x : std_logic_vector) return int816_t;
subtype uint817_t is unsigned(816 downto 0);
constant uint817_t_SLV_LEN : integer := 817;
function uint817_t_to_slv(x : uint817_t) return std_logic_vector;
function slv_to_uint817_t(x : std_logic_vector) return uint817_t;
subtype int817_t is signed(816 downto 0);
constant int817_t_SLV_LEN : integer := 817;
function int817_t_to_slv(x : int817_t) return std_logic_vector;
function slv_to_int817_t(x : std_logic_vector) return int817_t;
subtype uint818_t is unsigned(817 downto 0);
constant uint818_t_SLV_LEN : integer := 818;
function uint818_t_to_slv(x : uint818_t) return std_logic_vector;
function slv_to_uint818_t(x : std_logic_vector) return uint818_t;
subtype int818_t is signed(817 downto 0);
constant int818_t_SLV_LEN : integer := 818;
function int818_t_to_slv(x : int818_t) return std_logic_vector;
function slv_to_int818_t(x : std_logic_vector) return int818_t;
subtype uint819_t is unsigned(818 downto 0);
constant uint819_t_SLV_LEN : integer := 819;
function uint819_t_to_slv(x : uint819_t) return std_logic_vector;
function slv_to_uint819_t(x : std_logic_vector) return uint819_t;
subtype int819_t is signed(818 downto 0);
constant int819_t_SLV_LEN : integer := 819;
function int819_t_to_slv(x : int819_t) return std_logic_vector;
function slv_to_int819_t(x : std_logic_vector) return int819_t;
subtype uint820_t is unsigned(819 downto 0);
constant uint820_t_SLV_LEN : integer := 820;
function uint820_t_to_slv(x : uint820_t) return std_logic_vector;
function slv_to_uint820_t(x : std_logic_vector) return uint820_t;
subtype int820_t is signed(819 downto 0);
constant int820_t_SLV_LEN : integer := 820;
function int820_t_to_slv(x : int820_t) return std_logic_vector;
function slv_to_int820_t(x : std_logic_vector) return int820_t;
subtype uint821_t is unsigned(820 downto 0);
constant uint821_t_SLV_LEN : integer := 821;
function uint821_t_to_slv(x : uint821_t) return std_logic_vector;
function slv_to_uint821_t(x : std_logic_vector) return uint821_t;
subtype int821_t is signed(820 downto 0);
constant int821_t_SLV_LEN : integer := 821;
function int821_t_to_slv(x : int821_t) return std_logic_vector;
function slv_to_int821_t(x : std_logic_vector) return int821_t;
subtype uint822_t is unsigned(821 downto 0);
constant uint822_t_SLV_LEN : integer := 822;
function uint822_t_to_slv(x : uint822_t) return std_logic_vector;
function slv_to_uint822_t(x : std_logic_vector) return uint822_t;
subtype int822_t is signed(821 downto 0);
constant int822_t_SLV_LEN : integer := 822;
function int822_t_to_slv(x : int822_t) return std_logic_vector;
function slv_to_int822_t(x : std_logic_vector) return int822_t;
subtype uint823_t is unsigned(822 downto 0);
constant uint823_t_SLV_LEN : integer := 823;
function uint823_t_to_slv(x : uint823_t) return std_logic_vector;
function slv_to_uint823_t(x : std_logic_vector) return uint823_t;
subtype int823_t is signed(822 downto 0);
constant int823_t_SLV_LEN : integer := 823;
function int823_t_to_slv(x : int823_t) return std_logic_vector;
function slv_to_int823_t(x : std_logic_vector) return int823_t;
subtype uint824_t is unsigned(823 downto 0);
constant uint824_t_SLV_LEN : integer := 824;
function uint824_t_to_slv(x : uint824_t) return std_logic_vector;
function slv_to_uint824_t(x : std_logic_vector) return uint824_t;
subtype int824_t is signed(823 downto 0);
constant int824_t_SLV_LEN : integer := 824;
function int824_t_to_slv(x : int824_t) return std_logic_vector;
function slv_to_int824_t(x : std_logic_vector) return int824_t;
subtype uint825_t is unsigned(824 downto 0);
constant uint825_t_SLV_LEN : integer := 825;
function uint825_t_to_slv(x : uint825_t) return std_logic_vector;
function slv_to_uint825_t(x : std_logic_vector) return uint825_t;
subtype int825_t is signed(824 downto 0);
constant int825_t_SLV_LEN : integer := 825;
function int825_t_to_slv(x : int825_t) return std_logic_vector;
function slv_to_int825_t(x : std_logic_vector) return int825_t;
subtype uint826_t is unsigned(825 downto 0);
constant uint826_t_SLV_LEN : integer := 826;
function uint826_t_to_slv(x : uint826_t) return std_logic_vector;
function slv_to_uint826_t(x : std_logic_vector) return uint826_t;
subtype int826_t is signed(825 downto 0);
constant int826_t_SLV_LEN : integer := 826;
function int826_t_to_slv(x : int826_t) return std_logic_vector;
function slv_to_int826_t(x : std_logic_vector) return int826_t;
subtype uint827_t is unsigned(826 downto 0);
constant uint827_t_SLV_LEN : integer := 827;
function uint827_t_to_slv(x : uint827_t) return std_logic_vector;
function slv_to_uint827_t(x : std_logic_vector) return uint827_t;
subtype int827_t is signed(826 downto 0);
constant int827_t_SLV_LEN : integer := 827;
function int827_t_to_slv(x : int827_t) return std_logic_vector;
function slv_to_int827_t(x : std_logic_vector) return int827_t;
subtype uint828_t is unsigned(827 downto 0);
constant uint828_t_SLV_LEN : integer := 828;
function uint828_t_to_slv(x : uint828_t) return std_logic_vector;
function slv_to_uint828_t(x : std_logic_vector) return uint828_t;
subtype int828_t is signed(827 downto 0);
constant int828_t_SLV_LEN : integer := 828;
function int828_t_to_slv(x : int828_t) return std_logic_vector;
function slv_to_int828_t(x : std_logic_vector) return int828_t;
subtype uint829_t is unsigned(828 downto 0);
constant uint829_t_SLV_LEN : integer := 829;
function uint829_t_to_slv(x : uint829_t) return std_logic_vector;
function slv_to_uint829_t(x : std_logic_vector) return uint829_t;
subtype int829_t is signed(828 downto 0);
constant int829_t_SLV_LEN : integer := 829;
function int829_t_to_slv(x : int829_t) return std_logic_vector;
function slv_to_int829_t(x : std_logic_vector) return int829_t;
subtype uint830_t is unsigned(829 downto 0);
constant uint830_t_SLV_LEN : integer := 830;
function uint830_t_to_slv(x : uint830_t) return std_logic_vector;
function slv_to_uint830_t(x : std_logic_vector) return uint830_t;
subtype int830_t is signed(829 downto 0);
constant int830_t_SLV_LEN : integer := 830;
function int830_t_to_slv(x : int830_t) return std_logic_vector;
function slv_to_int830_t(x : std_logic_vector) return int830_t;
subtype uint831_t is unsigned(830 downto 0);
constant uint831_t_SLV_LEN : integer := 831;
function uint831_t_to_slv(x : uint831_t) return std_logic_vector;
function slv_to_uint831_t(x : std_logic_vector) return uint831_t;
subtype int831_t is signed(830 downto 0);
constant int831_t_SLV_LEN : integer := 831;
function int831_t_to_slv(x : int831_t) return std_logic_vector;
function slv_to_int831_t(x : std_logic_vector) return int831_t;
subtype uint832_t is unsigned(831 downto 0);
constant uint832_t_SLV_LEN : integer := 832;
function uint832_t_to_slv(x : uint832_t) return std_logic_vector;
function slv_to_uint832_t(x : std_logic_vector) return uint832_t;
subtype int832_t is signed(831 downto 0);
constant int832_t_SLV_LEN : integer := 832;
function int832_t_to_slv(x : int832_t) return std_logic_vector;
function slv_to_int832_t(x : std_logic_vector) return int832_t;
subtype uint833_t is unsigned(832 downto 0);
constant uint833_t_SLV_LEN : integer := 833;
function uint833_t_to_slv(x : uint833_t) return std_logic_vector;
function slv_to_uint833_t(x : std_logic_vector) return uint833_t;
subtype int833_t is signed(832 downto 0);
constant int833_t_SLV_LEN : integer := 833;
function int833_t_to_slv(x : int833_t) return std_logic_vector;
function slv_to_int833_t(x : std_logic_vector) return int833_t;
subtype uint834_t is unsigned(833 downto 0);
constant uint834_t_SLV_LEN : integer := 834;
function uint834_t_to_slv(x : uint834_t) return std_logic_vector;
function slv_to_uint834_t(x : std_logic_vector) return uint834_t;
subtype int834_t is signed(833 downto 0);
constant int834_t_SLV_LEN : integer := 834;
function int834_t_to_slv(x : int834_t) return std_logic_vector;
function slv_to_int834_t(x : std_logic_vector) return int834_t;
subtype uint835_t is unsigned(834 downto 0);
constant uint835_t_SLV_LEN : integer := 835;
function uint835_t_to_slv(x : uint835_t) return std_logic_vector;
function slv_to_uint835_t(x : std_logic_vector) return uint835_t;
subtype int835_t is signed(834 downto 0);
constant int835_t_SLV_LEN : integer := 835;
function int835_t_to_slv(x : int835_t) return std_logic_vector;
function slv_to_int835_t(x : std_logic_vector) return int835_t;
subtype uint836_t is unsigned(835 downto 0);
constant uint836_t_SLV_LEN : integer := 836;
function uint836_t_to_slv(x : uint836_t) return std_logic_vector;
function slv_to_uint836_t(x : std_logic_vector) return uint836_t;
subtype int836_t is signed(835 downto 0);
constant int836_t_SLV_LEN : integer := 836;
function int836_t_to_slv(x : int836_t) return std_logic_vector;
function slv_to_int836_t(x : std_logic_vector) return int836_t;
subtype uint837_t is unsigned(836 downto 0);
constant uint837_t_SLV_LEN : integer := 837;
function uint837_t_to_slv(x : uint837_t) return std_logic_vector;
function slv_to_uint837_t(x : std_logic_vector) return uint837_t;
subtype int837_t is signed(836 downto 0);
constant int837_t_SLV_LEN : integer := 837;
function int837_t_to_slv(x : int837_t) return std_logic_vector;
function slv_to_int837_t(x : std_logic_vector) return int837_t;
subtype uint838_t is unsigned(837 downto 0);
constant uint838_t_SLV_LEN : integer := 838;
function uint838_t_to_slv(x : uint838_t) return std_logic_vector;
function slv_to_uint838_t(x : std_logic_vector) return uint838_t;
subtype int838_t is signed(837 downto 0);
constant int838_t_SLV_LEN : integer := 838;
function int838_t_to_slv(x : int838_t) return std_logic_vector;
function slv_to_int838_t(x : std_logic_vector) return int838_t;
subtype uint839_t is unsigned(838 downto 0);
constant uint839_t_SLV_LEN : integer := 839;
function uint839_t_to_slv(x : uint839_t) return std_logic_vector;
function slv_to_uint839_t(x : std_logic_vector) return uint839_t;
subtype int839_t is signed(838 downto 0);
constant int839_t_SLV_LEN : integer := 839;
function int839_t_to_slv(x : int839_t) return std_logic_vector;
function slv_to_int839_t(x : std_logic_vector) return int839_t;
subtype uint840_t is unsigned(839 downto 0);
constant uint840_t_SLV_LEN : integer := 840;
function uint840_t_to_slv(x : uint840_t) return std_logic_vector;
function slv_to_uint840_t(x : std_logic_vector) return uint840_t;
subtype int840_t is signed(839 downto 0);
constant int840_t_SLV_LEN : integer := 840;
function int840_t_to_slv(x : int840_t) return std_logic_vector;
function slv_to_int840_t(x : std_logic_vector) return int840_t;
subtype uint841_t is unsigned(840 downto 0);
constant uint841_t_SLV_LEN : integer := 841;
function uint841_t_to_slv(x : uint841_t) return std_logic_vector;
function slv_to_uint841_t(x : std_logic_vector) return uint841_t;
subtype int841_t is signed(840 downto 0);
constant int841_t_SLV_LEN : integer := 841;
function int841_t_to_slv(x : int841_t) return std_logic_vector;
function slv_to_int841_t(x : std_logic_vector) return int841_t;
subtype uint842_t is unsigned(841 downto 0);
constant uint842_t_SLV_LEN : integer := 842;
function uint842_t_to_slv(x : uint842_t) return std_logic_vector;
function slv_to_uint842_t(x : std_logic_vector) return uint842_t;
subtype int842_t is signed(841 downto 0);
constant int842_t_SLV_LEN : integer := 842;
function int842_t_to_slv(x : int842_t) return std_logic_vector;
function slv_to_int842_t(x : std_logic_vector) return int842_t;
subtype uint843_t is unsigned(842 downto 0);
constant uint843_t_SLV_LEN : integer := 843;
function uint843_t_to_slv(x : uint843_t) return std_logic_vector;
function slv_to_uint843_t(x : std_logic_vector) return uint843_t;
subtype int843_t is signed(842 downto 0);
constant int843_t_SLV_LEN : integer := 843;
function int843_t_to_slv(x : int843_t) return std_logic_vector;
function slv_to_int843_t(x : std_logic_vector) return int843_t;
subtype uint844_t is unsigned(843 downto 0);
constant uint844_t_SLV_LEN : integer := 844;
function uint844_t_to_slv(x : uint844_t) return std_logic_vector;
function slv_to_uint844_t(x : std_logic_vector) return uint844_t;
subtype int844_t is signed(843 downto 0);
constant int844_t_SLV_LEN : integer := 844;
function int844_t_to_slv(x : int844_t) return std_logic_vector;
function slv_to_int844_t(x : std_logic_vector) return int844_t;
subtype uint845_t is unsigned(844 downto 0);
constant uint845_t_SLV_LEN : integer := 845;
function uint845_t_to_slv(x : uint845_t) return std_logic_vector;
function slv_to_uint845_t(x : std_logic_vector) return uint845_t;
subtype int845_t is signed(844 downto 0);
constant int845_t_SLV_LEN : integer := 845;
function int845_t_to_slv(x : int845_t) return std_logic_vector;
function slv_to_int845_t(x : std_logic_vector) return int845_t;
subtype uint846_t is unsigned(845 downto 0);
constant uint846_t_SLV_LEN : integer := 846;
function uint846_t_to_slv(x : uint846_t) return std_logic_vector;
function slv_to_uint846_t(x : std_logic_vector) return uint846_t;
subtype int846_t is signed(845 downto 0);
constant int846_t_SLV_LEN : integer := 846;
function int846_t_to_slv(x : int846_t) return std_logic_vector;
function slv_to_int846_t(x : std_logic_vector) return int846_t;
subtype uint847_t is unsigned(846 downto 0);
constant uint847_t_SLV_LEN : integer := 847;
function uint847_t_to_slv(x : uint847_t) return std_logic_vector;
function slv_to_uint847_t(x : std_logic_vector) return uint847_t;
subtype int847_t is signed(846 downto 0);
constant int847_t_SLV_LEN : integer := 847;
function int847_t_to_slv(x : int847_t) return std_logic_vector;
function slv_to_int847_t(x : std_logic_vector) return int847_t;
subtype uint848_t is unsigned(847 downto 0);
constant uint848_t_SLV_LEN : integer := 848;
function uint848_t_to_slv(x : uint848_t) return std_logic_vector;
function slv_to_uint848_t(x : std_logic_vector) return uint848_t;
subtype int848_t is signed(847 downto 0);
constant int848_t_SLV_LEN : integer := 848;
function int848_t_to_slv(x : int848_t) return std_logic_vector;
function slv_to_int848_t(x : std_logic_vector) return int848_t;
subtype uint849_t is unsigned(848 downto 0);
constant uint849_t_SLV_LEN : integer := 849;
function uint849_t_to_slv(x : uint849_t) return std_logic_vector;
function slv_to_uint849_t(x : std_logic_vector) return uint849_t;
subtype int849_t is signed(848 downto 0);
constant int849_t_SLV_LEN : integer := 849;
function int849_t_to_slv(x : int849_t) return std_logic_vector;
function slv_to_int849_t(x : std_logic_vector) return int849_t;
subtype uint850_t is unsigned(849 downto 0);
constant uint850_t_SLV_LEN : integer := 850;
function uint850_t_to_slv(x : uint850_t) return std_logic_vector;
function slv_to_uint850_t(x : std_logic_vector) return uint850_t;
subtype int850_t is signed(849 downto 0);
constant int850_t_SLV_LEN : integer := 850;
function int850_t_to_slv(x : int850_t) return std_logic_vector;
function slv_to_int850_t(x : std_logic_vector) return int850_t;
subtype uint851_t is unsigned(850 downto 0);
constant uint851_t_SLV_LEN : integer := 851;
function uint851_t_to_slv(x : uint851_t) return std_logic_vector;
function slv_to_uint851_t(x : std_logic_vector) return uint851_t;
subtype int851_t is signed(850 downto 0);
constant int851_t_SLV_LEN : integer := 851;
function int851_t_to_slv(x : int851_t) return std_logic_vector;
function slv_to_int851_t(x : std_logic_vector) return int851_t;
subtype uint852_t is unsigned(851 downto 0);
constant uint852_t_SLV_LEN : integer := 852;
function uint852_t_to_slv(x : uint852_t) return std_logic_vector;
function slv_to_uint852_t(x : std_logic_vector) return uint852_t;
subtype int852_t is signed(851 downto 0);
constant int852_t_SLV_LEN : integer := 852;
function int852_t_to_slv(x : int852_t) return std_logic_vector;
function slv_to_int852_t(x : std_logic_vector) return int852_t;
subtype uint853_t is unsigned(852 downto 0);
constant uint853_t_SLV_LEN : integer := 853;
function uint853_t_to_slv(x : uint853_t) return std_logic_vector;
function slv_to_uint853_t(x : std_logic_vector) return uint853_t;
subtype int853_t is signed(852 downto 0);
constant int853_t_SLV_LEN : integer := 853;
function int853_t_to_slv(x : int853_t) return std_logic_vector;
function slv_to_int853_t(x : std_logic_vector) return int853_t;
subtype uint854_t is unsigned(853 downto 0);
constant uint854_t_SLV_LEN : integer := 854;
function uint854_t_to_slv(x : uint854_t) return std_logic_vector;
function slv_to_uint854_t(x : std_logic_vector) return uint854_t;
subtype int854_t is signed(853 downto 0);
constant int854_t_SLV_LEN : integer := 854;
function int854_t_to_slv(x : int854_t) return std_logic_vector;
function slv_to_int854_t(x : std_logic_vector) return int854_t;
subtype uint855_t is unsigned(854 downto 0);
constant uint855_t_SLV_LEN : integer := 855;
function uint855_t_to_slv(x : uint855_t) return std_logic_vector;
function slv_to_uint855_t(x : std_logic_vector) return uint855_t;
subtype int855_t is signed(854 downto 0);
constant int855_t_SLV_LEN : integer := 855;
function int855_t_to_slv(x : int855_t) return std_logic_vector;
function slv_to_int855_t(x : std_logic_vector) return int855_t;
subtype uint856_t is unsigned(855 downto 0);
constant uint856_t_SLV_LEN : integer := 856;
function uint856_t_to_slv(x : uint856_t) return std_logic_vector;
function slv_to_uint856_t(x : std_logic_vector) return uint856_t;
subtype int856_t is signed(855 downto 0);
constant int856_t_SLV_LEN : integer := 856;
function int856_t_to_slv(x : int856_t) return std_logic_vector;
function slv_to_int856_t(x : std_logic_vector) return int856_t;
subtype uint857_t is unsigned(856 downto 0);
constant uint857_t_SLV_LEN : integer := 857;
function uint857_t_to_slv(x : uint857_t) return std_logic_vector;
function slv_to_uint857_t(x : std_logic_vector) return uint857_t;
subtype int857_t is signed(856 downto 0);
constant int857_t_SLV_LEN : integer := 857;
function int857_t_to_slv(x : int857_t) return std_logic_vector;
function slv_to_int857_t(x : std_logic_vector) return int857_t;
subtype uint858_t is unsigned(857 downto 0);
constant uint858_t_SLV_LEN : integer := 858;
function uint858_t_to_slv(x : uint858_t) return std_logic_vector;
function slv_to_uint858_t(x : std_logic_vector) return uint858_t;
subtype int858_t is signed(857 downto 0);
constant int858_t_SLV_LEN : integer := 858;
function int858_t_to_slv(x : int858_t) return std_logic_vector;
function slv_to_int858_t(x : std_logic_vector) return int858_t;
subtype uint859_t is unsigned(858 downto 0);
constant uint859_t_SLV_LEN : integer := 859;
function uint859_t_to_slv(x : uint859_t) return std_logic_vector;
function slv_to_uint859_t(x : std_logic_vector) return uint859_t;
subtype int859_t is signed(858 downto 0);
constant int859_t_SLV_LEN : integer := 859;
function int859_t_to_slv(x : int859_t) return std_logic_vector;
function slv_to_int859_t(x : std_logic_vector) return int859_t;
subtype uint860_t is unsigned(859 downto 0);
constant uint860_t_SLV_LEN : integer := 860;
function uint860_t_to_slv(x : uint860_t) return std_logic_vector;
function slv_to_uint860_t(x : std_logic_vector) return uint860_t;
subtype int860_t is signed(859 downto 0);
constant int860_t_SLV_LEN : integer := 860;
function int860_t_to_slv(x : int860_t) return std_logic_vector;
function slv_to_int860_t(x : std_logic_vector) return int860_t;
subtype uint861_t is unsigned(860 downto 0);
constant uint861_t_SLV_LEN : integer := 861;
function uint861_t_to_slv(x : uint861_t) return std_logic_vector;
function slv_to_uint861_t(x : std_logic_vector) return uint861_t;
subtype int861_t is signed(860 downto 0);
constant int861_t_SLV_LEN : integer := 861;
function int861_t_to_slv(x : int861_t) return std_logic_vector;
function slv_to_int861_t(x : std_logic_vector) return int861_t;
subtype uint862_t is unsigned(861 downto 0);
constant uint862_t_SLV_LEN : integer := 862;
function uint862_t_to_slv(x : uint862_t) return std_logic_vector;
function slv_to_uint862_t(x : std_logic_vector) return uint862_t;
subtype int862_t is signed(861 downto 0);
constant int862_t_SLV_LEN : integer := 862;
function int862_t_to_slv(x : int862_t) return std_logic_vector;
function slv_to_int862_t(x : std_logic_vector) return int862_t;
subtype uint863_t is unsigned(862 downto 0);
constant uint863_t_SLV_LEN : integer := 863;
function uint863_t_to_slv(x : uint863_t) return std_logic_vector;
function slv_to_uint863_t(x : std_logic_vector) return uint863_t;
subtype int863_t is signed(862 downto 0);
constant int863_t_SLV_LEN : integer := 863;
function int863_t_to_slv(x : int863_t) return std_logic_vector;
function slv_to_int863_t(x : std_logic_vector) return int863_t;
subtype uint864_t is unsigned(863 downto 0);
constant uint864_t_SLV_LEN : integer := 864;
function uint864_t_to_slv(x : uint864_t) return std_logic_vector;
function slv_to_uint864_t(x : std_logic_vector) return uint864_t;
subtype int864_t is signed(863 downto 0);
constant int864_t_SLV_LEN : integer := 864;
function int864_t_to_slv(x : int864_t) return std_logic_vector;
function slv_to_int864_t(x : std_logic_vector) return int864_t;
subtype uint865_t is unsigned(864 downto 0);
constant uint865_t_SLV_LEN : integer := 865;
function uint865_t_to_slv(x : uint865_t) return std_logic_vector;
function slv_to_uint865_t(x : std_logic_vector) return uint865_t;
subtype int865_t is signed(864 downto 0);
constant int865_t_SLV_LEN : integer := 865;
function int865_t_to_slv(x : int865_t) return std_logic_vector;
function slv_to_int865_t(x : std_logic_vector) return int865_t;
subtype uint866_t is unsigned(865 downto 0);
constant uint866_t_SLV_LEN : integer := 866;
function uint866_t_to_slv(x : uint866_t) return std_logic_vector;
function slv_to_uint866_t(x : std_logic_vector) return uint866_t;
subtype int866_t is signed(865 downto 0);
constant int866_t_SLV_LEN : integer := 866;
function int866_t_to_slv(x : int866_t) return std_logic_vector;
function slv_to_int866_t(x : std_logic_vector) return int866_t;
subtype uint867_t is unsigned(866 downto 0);
constant uint867_t_SLV_LEN : integer := 867;
function uint867_t_to_slv(x : uint867_t) return std_logic_vector;
function slv_to_uint867_t(x : std_logic_vector) return uint867_t;
subtype int867_t is signed(866 downto 0);
constant int867_t_SLV_LEN : integer := 867;
function int867_t_to_slv(x : int867_t) return std_logic_vector;
function slv_to_int867_t(x : std_logic_vector) return int867_t;
subtype uint868_t is unsigned(867 downto 0);
constant uint868_t_SLV_LEN : integer := 868;
function uint868_t_to_slv(x : uint868_t) return std_logic_vector;
function slv_to_uint868_t(x : std_logic_vector) return uint868_t;
subtype int868_t is signed(867 downto 0);
constant int868_t_SLV_LEN : integer := 868;
function int868_t_to_slv(x : int868_t) return std_logic_vector;
function slv_to_int868_t(x : std_logic_vector) return int868_t;
subtype uint869_t is unsigned(868 downto 0);
constant uint869_t_SLV_LEN : integer := 869;
function uint869_t_to_slv(x : uint869_t) return std_logic_vector;
function slv_to_uint869_t(x : std_logic_vector) return uint869_t;
subtype int869_t is signed(868 downto 0);
constant int869_t_SLV_LEN : integer := 869;
function int869_t_to_slv(x : int869_t) return std_logic_vector;
function slv_to_int869_t(x : std_logic_vector) return int869_t;
subtype uint870_t is unsigned(869 downto 0);
constant uint870_t_SLV_LEN : integer := 870;
function uint870_t_to_slv(x : uint870_t) return std_logic_vector;
function slv_to_uint870_t(x : std_logic_vector) return uint870_t;
subtype int870_t is signed(869 downto 0);
constant int870_t_SLV_LEN : integer := 870;
function int870_t_to_slv(x : int870_t) return std_logic_vector;
function slv_to_int870_t(x : std_logic_vector) return int870_t;
subtype uint871_t is unsigned(870 downto 0);
constant uint871_t_SLV_LEN : integer := 871;
function uint871_t_to_slv(x : uint871_t) return std_logic_vector;
function slv_to_uint871_t(x : std_logic_vector) return uint871_t;
subtype int871_t is signed(870 downto 0);
constant int871_t_SLV_LEN : integer := 871;
function int871_t_to_slv(x : int871_t) return std_logic_vector;
function slv_to_int871_t(x : std_logic_vector) return int871_t;
subtype uint872_t is unsigned(871 downto 0);
constant uint872_t_SLV_LEN : integer := 872;
function uint872_t_to_slv(x : uint872_t) return std_logic_vector;
function slv_to_uint872_t(x : std_logic_vector) return uint872_t;
subtype int872_t is signed(871 downto 0);
constant int872_t_SLV_LEN : integer := 872;
function int872_t_to_slv(x : int872_t) return std_logic_vector;
function slv_to_int872_t(x : std_logic_vector) return int872_t;
subtype uint873_t is unsigned(872 downto 0);
constant uint873_t_SLV_LEN : integer := 873;
function uint873_t_to_slv(x : uint873_t) return std_logic_vector;
function slv_to_uint873_t(x : std_logic_vector) return uint873_t;
subtype int873_t is signed(872 downto 0);
constant int873_t_SLV_LEN : integer := 873;
function int873_t_to_slv(x : int873_t) return std_logic_vector;
function slv_to_int873_t(x : std_logic_vector) return int873_t;
subtype uint874_t is unsigned(873 downto 0);
constant uint874_t_SLV_LEN : integer := 874;
function uint874_t_to_slv(x : uint874_t) return std_logic_vector;
function slv_to_uint874_t(x : std_logic_vector) return uint874_t;
subtype int874_t is signed(873 downto 0);
constant int874_t_SLV_LEN : integer := 874;
function int874_t_to_slv(x : int874_t) return std_logic_vector;
function slv_to_int874_t(x : std_logic_vector) return int874_t;
subtype uint875_t is unsigned(874 downto 0);
constant uint875_t_SLV_LEN : integer := 875;
function uint875_t_to_slv(x : uint875_t) return std_logic_vector;
function slv_to_uint875_t(x : std_logic_vector) return uint875_t;
subtype int875_t is signed(874 downto 0);
constant int875_t_SLV_LEN : integer := 875;
function int875_t_to_slv(x : int875_t) return std_logic_vector;
function slv_to_int875_t(x : std_logic_vector) return int875_t;
subtype uint876_t is unsigned(875 downto 0);
constant uint876_t_SLV_LEN : integer := 876;
function uint876_t_to_slv(x : uint876_t) return std_logic_vector;
function slv_to_uint876_t(x : std_logic_vector) return uint876_t;
subtype int876_t is signed(875 downto 0);
constant int876_t_SLV_LEN : integer := 876;
function int876_t_to_slv(x : int876_t) return std_logic_vector;
function slv_to_int876_t(x : std_logic_vector) return int876_t;
subtype uint877_t is unsigned(876 downto 0);
constant uint877_t_SLV_LEN : integer := 877;
function uint877_t_to_slv(x : uint877_t) return std_logic_vector;
function slv_to_uint877_t(x : std_logic_vector) return uint877_t;
subtype int877_t is signed(876 downto 0);
constant int877_t_SLV_LEN : integer := 877;
function int877_t_to_slv(x : int877_t) return std_logic_vector;
function slv_to_int877_t(x : std_logic_vector) return int877_t;
subtype uint878_t is unsigned(877 downto 0);
constant uint878_t_SLV_LEN : integer := 878;
function uint878_t_to_slv(x : uint878_t) return std_logic_vector;
function slv_to_uint878_t(x : std_logic_vector) return uint878_t;
subtype int878_t is signed(877 downto 0);
constant int878_t_SLV_LEN : integer := 878;
function int878_t_to_slv(x : int878_t) return std_logic_vector;
function slv_to_int878_t(x : std_logic_vector) return int878_t;
subtype uint879_t is unsigned(878 downto 0);
constant uint879_t_SLV_LEN : integer := 879;
function uint879_t_to_slv(x : uint879_t) return std_logic_vector;
function slv_to_uint879_t(x : std_logic_vector) return uint879_t;
subtype int879_t is signed(878 downto 0);
constant int879_t_SLV_LEN : integer := 879;
function int879_t_to_slv(x : int879_t) return std_logic_vector;
function slv_to_int879_t(x : std_logic_vector) return int879_t;
subtype uint880_t is unsigned(879 downto 0);
constant uint880_t_SLV_LEN : integer := 880;
function uint880_t_to_slv(x : uint880_t) return std_logic_vector;
function slv_to_uint880_t(x : std_logic_vector) return uint880_t;
subtype int880_t is signed(879 downto 0);
constant int880_t_SLV_LEN : integer := 880;
function int880_t_to_slv(x : int880_t) return std_logic_vector;
function slv_to_int880_t(x : std_logic_vector) return int880_t;
subtype uint881_t is unsigned(880 downto 0);
constant uint881_t_SLV_LEN : integer := 881;
function uint881_t_to_slv(x : uint881_t) return std_logic_vector;
function slv_to_uint881_t(x : std_logic_vector) return uint881_t;
subtype int881_t is signed(880 downto 0);
constant int881_t_SLV_LEN : integer := 881;
function int881_t_to_slv(x : int881_t) return std_logic_vector;
function slv_to_int881_t(x : std_logic_vector) return int881_t;
subtype uint882_t is unsigned(881 downto 0);
constant uint882_t_SLV_LEN : integer := 882;
function uint882_t_to_slv(x : uint882_t) return std_logic_vector;
function slv_to_uint882_t(x : std_logic_vector) return uint882_t;
subtype int882_t is signed(881 downto 0);
constant int882_t_SLV_LEN : integer := 882;
function int882_t_to_slv(x : int882_t) return std_logic_vector;
function slv_to_int882_t(x : std_logic_vector) return int882_t;
subtype uint883_t is unsigned(882 downto 0);
constant uint883_t_SLV_LEN : integer := 883;
function uint883_t_to_slv(x : uint883_t) return std_logic_vector;
function slv_to_uint883_t(x : std_logic_vector) return uint883_t;
subtype int883_t is signed(882 downto 0);
constant int883_t_SLV_LEN : integer := 883;
function int883_t_to_slv(x : int883_t) return std_logic_vector;
function slv_to_int883_t(x : std_logic_vector) return int883_t;
subtype uint884_t is unsigned(883 downto 0);
constant uint884_t_SLV_LEN : integer := 884;
function uint884_t_to_slv(x : uint884_t) return std_logic_vector;
function slv_to_uint884_t(x : std_logic_vector) return uint884_t;
subtype int884_t is signed(883 downto 0);
constant int884_t_SLV_LEN : integer := 884;
function int884_t_to_slv(x : int884_t) return std_logic_vector;
function slv_to_int884_t(x : std_logic_vector) return int884_t;
subtype uint885_t is unsigned(884 downto 0);
constant uint885_t_SLV_LEN : integer := 885;
function uint885_t_to_slv(x : uint885_t) return std_logic_vector;
function slv_to_uint885_t(x : std_logic_vector) return uint885_t;
subtype int885_t is signed(884 downto 0);
constant int885_t_SLV_LEN : integer := 885;
function int885_t_to_slv(x : int885_t) return std_logic_vector;
function slv_to_int885_t(x : std_logic_vector) return int885_t;
subtype uint886_t is unsigned(885 downto 0);
constant uint886_t_SLV_LEN : integer := 886;
function uint886_t_to_slv(x : uint886_t) return std_logic_vector;
function slv_to_uint886_t(x : std_logic_vector) return uint886_t;
subtype int886_t is signed(885 downto 0);
constant int886_t_SLV_LEN : integer := 886;
function int886_t_to_slv(x : int886_t) return std_logic_vector;
function slv_to_int886_t(x : std_logic_vector) return int886_t;
subtype uint887_t is unsigned(886 downto 0);
constant uint887_t_SLV_LEN : integer := 887;
function uint887_t_to_slv(x : uint887_t) return std_logic_vector;
function slv_to_uint887_t(x : std_logic_vector) return uint887_t;
subtype int887_t is signed(886 downto 0);
constant int887_t_SLV_LEN : integer := 887;
function int887_t_to_slv(x : int887_t) return std_logic_vector;
function slv_to_int887_t(x : std_logic_vector) return int887_t;
subtype uint888_t is unsigned(887 downto 0);
constant uint888_t_SLV_LEN : integer := 888;
function uint888_t_to_slv(x : uint888_t) return std_logic_vector;
function slv_to_uint888_t(x : std_logic_vector) return uint888_t;
subtype int888_t is signed(887 downto 0);
constant int888_t_SLV_LEN : integer := 888;
function int888_t_to_slv(x : int888_t) return std_logic_vector;
function slv_to_int888_t(x : std_logic_vector) return int888_t;
subtype uint889_t is unsigned(888 downto 0);
constant uint889_t_SLV_LEN : integer := 889;
function uint889_t_to_slv(x : uint889_t) return std_logic_vector;
function slv_to_uint889_t(x : std_logic_vector) return uint889_t;
subtype int889_t is signed(888 downto 0);
constant int889_t_SLV_LEN : integer := 889;
function int889_t_to_slv(x : int889_t) return std_logic_vector;
function slv_to_int889_t(x : std_logic_vector) return int889_t;
subtype uint890_t is unsigned(889 downto 0);
constant uint890_t_SLV_LEN : integer := 890;
function uint890_t_to_slv(x : uint890_t) return std_logic_vector;
function slv_to_uint890_t(x : std_logic_vector) return uint890_t;
subtype int890_t is signed(889 downto 0);
constant int890_t_SLV_LEN : integer := 890;
function int890_t_to_slv(x : int890_t) return std_logic_vector;
function slv_to_int890_t(x : std_logic_vector) return int890_t;
subtype uint891_t is unsigned(890 downto 0);
constant uint891_t_SLV_LEN : integer := 891;
function uint891_t_to_slv(x : uint891_t) return std_logic_vector;
function slv_to_uint891_t(x : std_logic_vector) return uint891_t;
subtype int891_t is signed(890 downto 0);
constant int891_t_SLV_LEN : integer := 891;
function int891_t_to_slv(x : int891_t) return std_logic_vector;
function slv_to_int891_t(x : std_logic_vector) return int891_t;
subtype uint892_t is unsigned(891 downto 0);
constant uint892_t_SLV_LEN : integer := 892;
function uint892_t_to_slv(x : uint892_t) return std_logic_vector;
function slv_to_uint892_t(x : std_logic_vector) return uint892_t;
subtype int892_t is signed(891 downto 0);
constant int892_t_SLV_LEN : integer := 892;
function int892_t_to_slv(x : int892_t) return std_logic_vector;
function slv_to_int892_t(x : std_logic_vector) return int892_t;
subtype uint893_t is unsigned(892 downto 0);
constant uint893_t_SLV_LEN : integer := 893;
function uint893_t_to_slv(x : uint893_t) return std_logic_vector;
function slv_to_uint893_t(x : std_logic_vector) return uint893_t;
subtype int893_t is signed(892 downto 0);
constant int893_t_SLV_LEN : integer := 893;
function int893_t_to_slv(x : int893_t) return std_logic_vector;
function slv_to_int893_t(x : std_logic_vector) return int893_t;
subtype uint894_t is unsigned(893 downto 0);
constant uint894_t_SLV_LEN : integer := 894;
function uint894_t_to_slv(x : uint894_t) return std_logic_vector;
function slv_to_uint894_t(x : std_logic_vector) return uint894_t;
subtype int894_t is signed(893 downto 0);
constant int894_t_SLV_LEN : integer := 894;
function int894_t_to_slv(x : int894_t) return std_logic_vector;
function slv_to_int894_t(x : std_logic_vector) return int894_t;
subtype uint895_t is unsigned(894 downto 0);
constant uint895_t_SLV_LEN : integer := 895;
function uint895_t_to_slv(x : uint895_t) return std_logic_vector;
function slv_to_uint895_t(x : std_logic_vector) return uint895_t;
subtype int895_t is signed(894 downto 0);
constant int895_t_SLV_LEN : integer := 895;
function int895_t_to_slv(x : int895_t) return std_logic_vector;
function slv_to_int895_t(x : std_logic_vector) return int895_t;
subtype uint896_t is unsigned(895 downto 0);
constant uint896_t_SLV_LEN : integer := 896;
function uint896_t_to_slv(x : uint896_t) return std_logic_vector;
function slv_to_uint896_t(x : std_logic_vector) return uint896_t;
subtype int896_t is signed(895 downto 0);
constant int896_t_SLV_LEN : integer := 896;
function int896_t_to_slv(x : int896_t) return std_logic_vector;
function slv_to_int896_t(x : std_logic_vector) return int896_t;
subtype uint897_t is unsigned(896 downto 0);
constant uint897_t_SLV_LEN : integer := 897;
function uint897_t_to_slv(x : uint897_t) return std_logic_vector;
function slv_to_uint897_t(x : std_logic_vector) return uint897_t;
subtype int897_t is signed(896 downto 0);
constant int897_t_SLV_LEN : integer := 897;
function int897_t_to_slv(x : int897_t) return std_logic_vector;
function slv_to_int897_t(x : std_logic_vector) return int897_t;
subtype uint898_t is unsigned(897 downto 0);
constant uint898_t_SLV_LEN : integer := 898;
function uint898_t_to_slv(x : uint898_t) return std_logic_vector;
function slv_to_uint898_t(x : std_logic_vector) return uint898_t;
subtype int898_t is signed(897 downto 0);
constant int898_t_SLV_LEN : integer := 898;
function int898_t_to_slv(x : int898_t) return std_logic_vector;
function slv_to_int898_t(x : std_logic_vector) return int898_t;
subtype uint899_t is unsigned(898 downto 0);
constant uint899_t_SLV_LEN : integer := 899;
function uint899_t_to_slv(x : uint899_t) return std_logic_vector;
function slv_to_uint899_t(x : std_logic_vector) return uint899_t;
subtype int899_t is signed(898 downto 0);
constant int899_t_SLV_LEN : integer := 899;
function int899_t_to_slv(x : int899_t) return std_logic_vector;
function slv_to_int899_t(x : std_logic_vector) return int899_t;
subtype uint900_t is unsigned(899 downto 0);
constant uint900_t_SLV_LEN : integer := 900;
function uint900_t_to_slv(x : uint900_t) return std_logic_vector;
function slv_to_uint900_t(x : std_logic_vector) return uint900_t;
subtype int900_t is signed(899 downto 0);
constant int900_t_SLV_LEN : integer := 900;
function int900_t_to_slv(x : int900_t) return std_logic_vector;
function slv_to_int900_t(x : std_logic_vector) return int900_t;
subtype uint901_t is unsigned(900 downto 0);
constant uint901_t_SLV_LEN : integer := 901;
function uint901_t_to_slv(x : uint901_t) return std_logic_vector;
function slv_to_uint901_t(x : std_logic_vector) return uint901_t;
subtype int901_t is signed(900 downto 0);
constant int901_t_SLV_LEN : integer := 901;
function int901_t_to_slv(x : int901_t) return std_logic_vector;
function slv_to_int901_t(x : std_logic_vector) return int901_t;
subtype uint902_t is unsigned(901 downto 0);
constant uint902_t_SLV_LEN : integer := 902;
function uint902_t_to_slv(x : uint902_t) return std_logic_vector;
function slv_to_uint902_t(x : std_logic_vector) return uint902_t;
subtype int902_t is signed(901 downto 0);
constant int902_t_SLV_LEN : integer := 902;
function int902_t_to_slv(x : int902_t) return std_logic_vector;
function slv_to_int902_t(x : std_logic_vector) return int902_t;
subtype uint903_t is unsigned(902 downto 0);
constant uint903_t_SLV_LEN : integer := 903;
function uint903_t_to_slv(x : uint903_t) return std_logic_vector;
function slv_to_uint903_t(x : std_logic_vector) return uint903_t;
subtype int903_t is signed(902 downto 0);
constant int903_t_SLV_LEN : integer := 903;
function int903_t_to_slv(x : int903_t) return std_logic_vector;
function slv_to_int903_t(x : std_logic_vector) return int903_t;
subtype uint904_t is unsigned(903 downto 0);
constant uint904_t_SLV_LEN : integer := 904;
function uint904_t_to_slv(x : uint904_t) return std_logic_vector;
function slv_to_uint904_t(x : std_logic_vector) return uint904_t;
subtype int904_t is signed(903 downto 0);
constant int904_t_SLV_LEN : integer := 904;
function int904_t_to_slv(x : int904_t) return std_logic_vector;
function slv_to_int904_t(x : std_logic_vector) return int904_t;
subtype uint905_t is unsigned(904 downto 0);
constant uint905_t_SLV_LEN : integer := 905;
function uint905_t_to_slv(x : uint905_t) return std_logic_vector;
function slv_to_uint905_t(x : std_logic_vector) return uint905_t;
subtype int905_t is signed(904 downto 0);
constant int905_t_SLV_LEN : integer := 905;
function int905_t_to_slv(x : int905_t) return std_logic_vector;
function slv_to_int905_t(x : std_logic_vector) return int905_t;
subtype uint906_t is unsigned(905 downto 0);
constant uint906_t_SLV_LEN : integer := 906;
function uint906_t_to_slv(x : uint906_t) return std_logic_vector;
function slv_to_uint906_t(x : std_logic_vector) return uint906_t;
subtype int906_t is signed(905 downto 0);
constant int906_t_SLV_LEN : integer := 906;
function int906_t_to_slv(x : int906_t) return std_logic_vector;
function slv_to_int906_t(x : std_logic_vector) return int906_t;
subtype uint907_t is unsigned(906 downto 0);
constant uint907_t_SLV_LEN : integer := 907;
function uint907_t_to_slv(x : uint907_t) return std_logic_vector;
function slv_to_uint907_t(x : std_logic_vector) return uint907_t;
subtype int907_t is signed(906 downto 0);
constant int907_t_SLV_LEN : integer := 907;
function int907_t_to_slv(x : int907_t) return std_logic_vector;
function slv_to_int907_t(x : std_logic_vector) return int907_t;
subtype uint908_t is unsigned(907 downto 0);
constant uint908_t_SLV_LEN : integer := 908;
function uint908_t_to_slv(x : uint908_t) return std_logic_vector;
function slv_to_uint908_t(x : std_logic_vector) return uint908_t;
subtype int908_t is signed(907 downto 0);
constant int908_t_SLV_LEN : integer := 908;
function int908_t_to_slv(x : int908_t) return std_logic_vector;
function slv_to_int908_t(x : std_logic_vector) return int908_t;
subtype uint909_t is unsigned(908 downto 0);
constant uint909_t_SLV_LEN : integer := 909;
function uint909_t_to_slv(x : uint909_t) return std_logic_vector;
function slv_to_uint909_t(x : std_logic_vector) return uint909_t;
subtype int909_t is signed(908 downto 0);
constant int909_t_SLV_LEN : integer := 909;
function int909_t_to_slv(x : int909_t) return std_logic_vector;
function slv_to_int909_t(x : std_logic_vector) return int909_t;
subtype uint910_t is unsigned(909 downto 0);
constant uint910_t_SLV_LEN : integer := 910;
function uint910_t_to_slv(x : uint910_t) return std_logic_vector;
function slv_to_uint910_t(x : std_logic_vector) return uint910_t;
subtype int910_t is signed(909 downto 0);
constant int910_t_SLV_LEN : integer := 910;
function int910_t_to_slv(x : int910_t) return std_logic_vector;
function slv_to_int910_t(x : std_logic_vector) return int910_t;
subtype uint911_t is unsigned(910 downto 0);
constant uint911_t_SLV_LEN : integer := 911;
function uint911_t_to_slv(x : uint911_t) return std_logic_vector;
function slv_to_uint911_t(x : std_logic_vector) return uint911_t;
subtype int911_t is signed(910 downto 0);
constant int911_t_SLV_LEN : integer := 911;
function int911_t_to_slv(x : int911_t) return std_logic_vector;
function slv_to_int911_t(x : std_logic_vector) return int911_t;
subtype uint912_t is unsigned(911 downto 0);
constant uint912_t_SLV_LEN : integer := 912;
function uint912_t_to_slv(x : uint912_t) return std_logic_vector;
function slv_to_uint912_t(x : std_logic_vector) return uint912_t;
subtype int912_t is signed(911 downto 0);
constant int912_t_SLV_LEN : integer := 912;
function int912_t_to_slv(x : int912_t) return std_logic_vector;
function slv_to_int912_t(x : std_logic_vector) return int912_t;
subtype uint913_t is unsigned(912 downto 0);
constant uint913_t_SLV_LEN : integer := 913;
function uint913_t_to_slv(x : uint913_t) return std_logic_vector;
function slv_to_uint913_t(x : std_logic_vector) return uint913_t;
subtype int913_t is signed(912 downto 0);
constant int913_t_SLV_LEN : integer := 913;
function int913_t_to_slv(x : int913_t) return std_logic_vector;
function slv_to_int913_t(x : std_logic_vector) return int913_t;
subtype uint914_t is unsigned(913 downto 0);
constant uint914_t_SLV_LEN : integer := 914;
function uint914_t_to_slv(x : uint914_t) return std_logic_vector;
function slv_to_uint914_t(x : std_logic_vector) return uint914_t;
subtype int914_t is signed(913 downto 0);
constant int914_t_SLV_LEN : integer := 914;
function int914_t_to_slv(x : int914_t) return std_logic_vector;
function slv_to_int914_t(x : std_logic_vector) return int914_t;
subtype uint915_t is unsigned(914 downto 0);
constant uint915_t_SLV_LEN : integer := 915;
function uint915_t_to_slv(x : uint915_t) return std_logic_vector;
function slv_to_uint915_t(x : std_logic_vector) return uint915_t;
subtype int915_t is signed(914 downto 0);
constant int915_t_SLV_LEN : integer := 915;
function int915_t_to_slv(x : int915_t) return std_logic_vector;
function slv_to_int915_t(x : std_logic_vector) return int915_t;
subtype uint916_t is unsigned(915 downto 0);
constant uint916_t_SLV_LEN : integer := 916;
function uint916_t_to_slv(x : uint916_t) return std_logic_vector;
function slv_to_uint916_t(x : std_logic_vector) return uint916_t;
subtype int916_t is signed(915 downto 0);
constant int916_t_SLV_LEN : integer := 916;
function int916_t_to_slv(x : int916_t) return std_logic_vector;
function slv_to_int916_t(x : std_logic_vector) return int916_t;
subtype uint917_t is unsigned(916 downto 0);
constant uint917_t_SLV_LEN : integer := 917;
function uint917_t_to_slv(x : uint917_t) return std_logic_vector;
function slv_to_uint917_t(x : std_logic_vector) return uint917_t;
subtype int917_t is signed(916 downto 0);
constant int917_t_SLV_LEN : integer := 917;
function int917_t_to_slv(x : int917_t) return std_logic_vector;
function slv_to_int917_t(x : std_logic_vector) return int917_t;
subtype uint918_t is unsigned(917 downto 0);
constant uint918_t_SLV_LEN : integer := 918;
function uint918_t_to_slv(x : uint918_t) return std_logic_vector;
function slv_to_uint918_t(x : std_logic_vector) return uint918_t;
subtype int918_t is signed(917 downto 0);
constant int918_t_SLV_LEN : integer := 918;
function int918_t_to_slv(x : int918_t) return std_logic_vector;
function slv_to_int918_t(x : std_logic_vector) return int918_t;
subtype uint919_t is unsigned(918 downto 0);
constant uint919_t_SLV_LEN : integer := 919;
function uint919_t_to_slv(x : uint919_t) return std_logic_vector;
function slv_to_uint919_t(x : std_logic_vector) return uint919_t;
subtype int919_t is signed(918 downto 0);
constant int919_t_SLV_LEN : integer := 919;
function int919_t_to_slv(x : int919_t) return std_logic_vector;
function slv_to_int919_t(x : std_logic_vector) return int919_t;
subtype uint920_t is unsigned(919 downto 0);
constant uint920_t_SLV_LEN : integer := 920;
function uint920_t_to_slv(x : uint920_t) return std_logic_vector;
function slv_to_uint920_t(x : std_logic_vector) return uint920_t;
subtype int920_t is signed(919 downto 0);
constant int920_t_SLV_LEN : integer := 920;
function int920_t_to_slv(x : int920_t) return std_logic_vector;
function slv_to_int920_t(x : std_logic_vector) return int920_t;
subtype uint921_t is unsigned(920 downto 0);
constant uint921_t_SLV_LEN : integer := 921;
function uint921_t_to_slv(x : uint921_t) return std_logic_vector;
function slv_to_uint921_t(x : std_logic_vector) return uint921_t;
subtype int921_t is signed(920 downto 0);
constant int921_t_SLV_LEN : integer := 921;
function int921_t_to_slv(x : int921_t) return std_logic_vector;
function slv_to_int921_t(x : std_logic_vector) return int921_t;
subtype uint922_t is unsigned(921 downto 0);
constant uint922_t_SLV_LEN : integer := 922;
function uint922_t_to_slv(x : uint922_t) return std_logic_vector;
function slv_to_uint922_t(x : std_logic_vector) return uint922_t;
subtype int922_t is signed(921 downto 0);
constant int922_t_SLV_LEN : integer := 922;
function int922_t_to_slv(x : int922_t) return std_logic_vector;
function slv_to_int922_t(x : std_logic_vector) return int922_t;
subtype uint923_t is unsigned(922 downto 0);
constant uint923_t_SLV_LEN : integer := 923;
function uint923_t_to_slv(x : uint923_t) return std_logic_vector;
function slv_to_uint923_t(x : std_logic_vector) return uint923_t;
subtype int923_t is signed(922 downto 0);
constant int923_t_SLV_LEN : integer := 923;
function int923_t_to_slv(x : int923_t) return std_logic_vector;
function slv_to_int923_t(x : std_logic_vector) return int923_t;
subtype uint924_t is unsigned(923 downto 0);
constant uint924_t_SLV_LEN : integer := 924;
function uint924_t_to_slv(x : uint924_t) return std_logic_vector;
function slv_to_uint924_t(x : std_logic_vector) return uint924_t;
subtype int924_t is signed(923 downto 0);
constant int924_t_SLV_LEN : integer := 924;
function int924_t_to_slv(x : int924_t) return std_logic_vector;
function slv_to_int924_t(x : std_logic_vector) return int924_t;
subtype uint925_t is unsigned(924 downto 0);
constant uint925_t_SLV_LEN : integer := 925;
function uint925_t_to_slv(x : uint925_t) return std_logic_vector;
function slv_to_uint925_t(x : std_logic_vector) return uint925_t;
subtype int925_t is signed(924 downto 0);
constant int925_t_SLV_LEN : integer := 925;
function int925_t_to_slv(x : int925_t) return std_logic_vector;
function slv_to_int925_t(x : std_logic_vector) return int925_t;
subtype uint926_t is unsigned(925 downto 0);
constant uint926_t_SLV_LEN : integer := 926;
function uint926_t_to_slv(x : uint926_t) return std_logic_vector;
function slv_to_uint926_t(x : std_logic_vector) return uint926_t;
subtype int926_t is signed(925 downto 0);
constant int926_t_SLV_LEN : integer := 926;
function int926_t_to_slv(x : int926_t) return std_logic_vector;
function slv_to_int926_t(x : std_logic_vector) return int926_t;
subtype uint927_t is unsigned(926 downto 0);
constant uint927_t_SLV_LEN : integer := 927;
function uint927_t_to_slv(x : uint927_t) return std_logic_vector;
function slv_to_uint927_t(x : std_logic_vector) return uint927_t;
subtype int927_t is signed(926 downto 0);
constant int927_t_SLV_LEN : integer := 927;
function int927_t_to_slv(x : int927_t) return std_logic_vector;
function slv_to_int927_t(x : std_logic_vector) return int927_t;
subtype uint928_t is unsigned(927 downto 0);
constant uint928_t_SLV_LEN : integer := 928;
function uint928_t_to_slv(x : uint928_t) return std_logic_vector;
function slv_to_uint928_t(x : std_logic_vector) return uint928_t;
subtype int928_t is signed(927 downto 0);
constant int928_t_SLV_LEN : integer := 928;
function int928_t_to_slv(x : int928_t) return std_logic_vector;
function slv_to_int928_t(x : std_logic_vector) return int928_t;
subtype uint929_t is unsigned(928 downto 0);
constant uint929_t_SLV_LEN : integer := 929;
function uint929_t_to_slv(x : uint929_t) return std_logic_vector;
function slv_to_uint929_t(x : std_logic_vector) return uint929_t;
subtype int929_t is signed(928 downto 0);
constant int929_t_SLV_LEN : integer := 929;
function int929_t_to_slv(x : int929_t) return std_logic_vector;
function slv_to_int929_t(x : std_logic_vector) return int929_t;
subtype uint930_t is unsigned(929 downto 0);
constant uint930_t_SLV_LEN : integer := 930;
function uint930_t_to_slv(x : uint930_t) return std_logic_vector;
function slv_to_uint930_t(x : std_logic_vector) return uint930_t;
subtype int930_t is signed(929 downto 0);
constant int930_t_SLV_LEN : integer := 930;
function int930_t_to_slv(x : int930_t) return std_logic_vector;
function slv_to_int930_t(x : std_logic_vector) return int930_t;
subtype uint931_t is unsigned(930 downto 0);
constant uint931_t_SLV_LEN : integer := 931;
function uint931_t_to_slv(x : uint931_t) return std_logic_vector;
function slv_to_uint931_t(x : std_logic_vector) return uint931_t;
subtype int931_t is signed(930 downto 0);
constant int931_t_SLV_LEN : integer := 931;
function int931_t_to_slv(x : int931_t) return std_logic_vector;
function slv_to_int931_t(x : std_logic_vector) return int931_t;
subtype uint932_t is unsigned(931 downto 0);
constant uint932_t_SLV_LEN : integer := 932;
function uint932_t_to_slv(x : uint932_t) return std_logic_vector;
function slv_to_uint932_t(x : std_logic_vector) return uint932_t;
subtype int932_t is signed(931 downto 0);
constant int932_t_SLV_LEN : integer := 932;
function int932_t_to_slv(x : int932_t) return std_logic_vector;
function slv_to_int932_t(x : std_logic_vector) return int932_t;
subtype uint933_t is unsigned(932 downto 0);
constant uint933_t_SLV_LEN : integer := 933;
function uint933_t_to_slv(x : uint933_t) return std_logic_vector;
function slv_to_uint933_t(x : std_logic_vector) return uint933_t;
subtype int933_t is signed(932 downto 0);
constant int933_t_SLV_LEN : integer := 933;
function int933_t_to_slv(x : int933_t) return std_logic_vector;
function slv_to_int933_t(x : std_logic_vector) return int933_t;
subtype uint934_t is unsigned(933 downto 0);
constant uint934_t_SLV_LEN : integer := 934;
function uint934_t_to_slv(x : uint934_t) return std_logic_vector;
function slv_to_uint934_t(x : std_logic_vector) return uint934_t;
subtype int934_t is signed(933 downto 0);
constant int934_t_SLV_LEN : integer := 934;
function int934_t_to_slv(x : int934_t) return std_logic_vector;
function slv_to_int934_t(x : std_logic_vector) return int934_t;
subtype uint935_t is unsigned(934 downto 0);
constant uint935_t_SLV_LEN : integer := 935;
function uint935_t_to_slv(x : uint935_t) return std_logic_vector;
function slv_to_uint935_t(x : std_logic_vector) return uint935_t;
subtype int935_t is signed(934 downto 0);
constant int935_t_SLV_LEN : integer := 935;
function int935_t_to_slv(x : int935_t) return std_logic_vector;
function slv_to_int935_t(x : std_logic_vector) return int935_t;
subtype uint936_t is unsigned(935 downto 0);
constant uint936_t_SLV_LEN : integer := 936;
function uint936_t_to_slv(x : uint936_t) return std_logic_vector;
function slv_to_uint936_t(x : std_logic_vector) return uint936_t;
subtype int936_t is signed(935 downto 0);
constant int936_t_SLV_LEN : integer := 936;
function int936_t_to_slv(x : int936_t) return std_logic_vector;
function slv_to_int936_t(x : std_logic_vector) return int936_t;
subtype uint937_t is unsigned(936 downto 0);
constant uint937_t_SLV_LEN : integer := 937;
function uint937_t_to_slv(x : uint937_t) return std_logic_vector;
function slv_to_uint937_t(x : std_logic_vector) return uint937_t;
subtype int937_t is signed(936 downto 0);
constant int937_t_SLV_LEN : integer := 937;
function int937_t_to_slv(x : int937_t) return std_logic_vector;
function slv_to_int937_t(x : std_logic_vector) return int937_t;
subtype uint938_t is unsigned(937 downto 0);
constant uint938_t_SLV_LEN : integer := 938;
function uint938_t_to_slv(x : uint938_t) return std_logic_vector;
function slv_to_uint938_t(x : std_logic_vector) return uint938_t;
subtype int938_t is signed(937 downto 0);
constant int938_t_SLV_LEN : integer := 938;
function int938_t_to_slv(x : int938_t) return std_logic_vector;
function slv_to_int938_t(x : std_logic_vector) return int938_t;
subtype uint939_t is unsigned(938 downto 0);
constant uint939_t_SLV_LEN : integer := 939;
function uint939_t_to_slv(x : uint939_t) return std_logic_vector;
function slv_to_uint939_t(x : std_logic_vector) return uint939_t;
subtype int939_t is signed(938 downto 0);
constant int939_t_SLV_LEN : integer := 939;
function int939_t_to_slv(x : int939_t) return std_logic_vector;
function slv_to_int939_t(x : std_logic_vector) return int939_t;
subtype uint940_t is unsigned(939 downto 0);
constant uint940_t_SLV_LEN : integer := 940;
function uint940_t_to_slv(x : uint940_t) return std_logic_vector;
function slv_to_uint940_t(x : std_logic_vector) return uint940_t;
subtype int940_t is signed(939 downto 0);
constant int940_t_SLV_LEN : integer := 940;
function int940_t_to_slv(x : int940_t) return std_logic_vector;
function slv_to_int940_t(x : std_logic_vector) return int940_t;
subtype uint941_t is unsigned(940 downto 0);
constant uint941_t_SLV_LEN : integer := 941;
function uint941_t_to_slv(x : uint941_t) return std_logic_vector;
function slv_to_uint941_t(x : std_logic_vector) return uint941_t;
subtype int941_t is signed(940 downto 0);
constant int941_t_SLV_LEN : integer := 941;
function int941_t_to_slv(x : int941_t) return std_logic_vector;
function slv_to_int941_t(x : std_logic_vector) return int941_t;
subtype uint942_t is unsigned(941 downto 0);
constant uint942_t_SLV_LEN : integer := 942;
function uint942_t_to_slv(x : uint942_t) return std_logic_vector;
function slv_to_uint942_t(x : std_logic_vector) return uint942_t;
subtype int942_t is signed(941 downto 0);
constant int942_t_SLV_LEN : integer := 942;
function int942_t_to_slv(x : int942_t) return std_logic_vector;
function slv_to_int942_t(x : std_logic_vector) return int942_t;
subtype uint943_t is unsigned(942 downto 0);
constant uint943_t_SLV_LEN : integer := 943;
function uint943_t_to_slv(x : uint943_t) return std_logic_vector;
function slv_to_uint943_t(x : std_logic_vector) return uint943_t;
subtype int943_t is signed(942 downto 0);
constant int943_t_SLV_LEN : integer := 943;
function int943_t_to_slv(x : int943_t) return std_logic_vector;
function slv_to_int943_t(x : std_logic_vector) return int943_t;
subtype uint944_t is unsigned(943 downto 0);
constant uint944_t_SLV_LEN : integer := 944;
function uint944_t_to_slv(x : uint944_t) return std_logic_vector;
function slv_to_uint944_t(x : std_logic_vector) return uint944_t;
subtype int944_t is signed(943 downto 0);
constant int944_t_SLV_LEN : integer := 944;
function int944_t_to_slv(x : int944_t) return std_logic_vector;
function slv_to_int944_t(x : std_logic_vector) return int944_t;
subtype uint945_t is unsigned(944 downto 0);
constant uint945_t_SLV_LEN : integer := 945;
function uint945_t_to_slv(x : uint945_t) return std_logic_vector;
function slv_to_uint945_t(x : std_logic_vector) return uint945_t;
subtype int945_t is signed(944 downto 0);
constant int945_t_SLV_LEN : integer := 945;
function int945_t_to_slv(x : int945_t) return std_logic_vector;
function slv_to_int945_t(x : std_logic_vector) return int945_t;
subtype uint946_t is unsigned(945 downto 0);
constant uint946_t_SLV_LEN : integer := 946;
function uint946_t_to_slv(x : uint946_t) return std_logic_vector;
function slv_to_uint946_t(x : std_logic_vector) return uint946_t;
subtype int946_t is signed(945 downto 0);
constant int946_t_SLV_LEN : integer := 946;
function int946_t_to_slv(x : int946_t) return std_logic_vector;
function slv_to_int946_t(x : std_logic_vector) return int946_t;
subtype uint947_t is unsigned(946 downto 0);
constant uint947_t_SLV_LEN : integer := 947;
function uint947_t_to_slv(x : uint947_t) return std_logic_vector;
function slv_to_uint947_t(x : std_logic_vector) return uint947_t;
subtype int947_t is signed(946 downto 0);
constant int947_t_SLV_LEN : integer := 947;
function int947_t_to_slv(x : int947_t) return std_logic_vector;
function slv_to_int947_t(x : std_logic_vector) return int947_t;
subtype uint948_t is unsigned(947 downto 0);
constant uint948_t_SLV_LEN : integer := 948;
function uint948_t_to_slv(x : uint948_t) return std_logic_vector;
function slv_to_uint948_t(x : std_logic_vector) return uint948_t;
subtype int948_t is signed(947 downto 0);
constant int948_t_SLV_LEN : integer := 948;
function int948_t_to_slv(x : int948_t) return std_logic_vector;
function slv_to_int948_t(x : std_logic_vector) return int948_t;
subtype uint949_t is unsigned(948 downto 0);
constant uint949_t_SLV_LEN : integer := 949;
function uint949_t_to_slv(x : uint949_t) return std_logic_vector;
function slv_to_uint949_t(x : std_logic_vector) return uint949_t;
subtype int949_t is signed(948 downto 0);
constant int949_t_SLV_LEN : integer := 949;
function int949_t_to_slv(x : int949_t) return std_logic_vector;
function slv_to_int949_t(x : std_logic_vector) return int949_t;
subtype uint950_t is unsigned(949 downto 0);
constant uint950_t_SLV_LEN : integer := 950;
function uint950_t_to_slv(x : uint950_t) return std_logic_vector;
function slv_to_uint950_t(x : std_logic_vector) return uint950_t;
subtype int950_t is signed(949 downto 0);
constant int950_t_SLV_LEN : integer := 950;
function int950_t_to_slv(x : int950_t) return std_logic_vector;
function slv_to_int950_t(x : std_logic_vector) return int950_t;
subtype uint951_t is unsigned(950 downto 0);
constant uint951_t_SLV_LEN : integer := 951;
function uint951_t_to_slv(x : uint951_t) return std_logic_vector;
function slv_to_uint951_t(x : std_logic_vector) return uint951_t;
subtype int951_t is signed(950 downto 0);
constant int951_t_SLV_LEN : integer := 951;
function int951_t_to_slv(x : int951_t) return std_logic_vector;
function slv_to_int951_t(x : std_logic_vector) return int951_t;
subtype uint952_t is unsigned(951 downto 0);
constant uint952_t_SLV_LEN : integer := 952;
function uint952_t_to_slv(x : uint952_t) return std_logic_vector;
function slv_to_uint952_t(x : std_logic_vector) return uint952_t;
subtype int952_t is signed(951 downto 0);
constant int952_t_SLV_LEN : integer := 952;
function int952_t_to_slv(x : int952_t) return std_logic_vector;
function slv_to_int952_t(x : std_logic_vector) return int952_t;
subtype uint953_t is unsigned(952 downto 0);
constant uint953_t_SLV_LEN : integer := 953;
function uint953_t_to_slv(x : uint953_t) return std_logic_vector;
function slv_to_uint953_t(x : std_logic_vector) return uint953_t;
subtype int953_t is signed(952 downto 0);
constant int953_t_SLV_LEN : integer := 953;
function int953_t_to_slv(x : int953_t) return std_logic_vector;
function slv_to_int953_t(x : std_logic_vector) return int953_t;
subtype uint954_t is unsigned(953 downto 0);
constant uint954_t_SLV_LEN : integer := 954;
function uint954_t_to_slv(x : uint954_t) return std_logic_vector;
function slv_to_uint954_t(x : std_logic_vector) return uint954_t;
subtype int954_t is signed(953 downto 0);
constant int954_t_SLV_LEN : integer := 954;
function int954_t_to_slv(x : int954_t) return std_logic_vector;
function slv_to_int954_t(x : std_logic_vector) return int954_t;
subtype uint955_t is unsigned(954 downto 0);
constant uint955_t_SLV_LEN : integer := 955;
function uint955_t_to_slv(x : uint955_t) return std_logic_vector;
function slv_to_uint955_t(x : std_logic_vector) return uint955_t;
subtype int955_t is signed(954 downto 0);
constant int955_t_SLV_LEN : integer := 955;
function int955_t_to_slv(x : int955_t) return std_logic_vector;
function slv_to_int955_t(x : std_logic_vector) return int955_t;
subtype uint956_t is unsigned(955 downto 0);
constant uint956_t_SLV_LEN : integer := 956;
function uint956_t_to_slv(x : uint956_t) return std_logic_vector;
function slv_to_uint956_t(x : std_logic_vector) return uint956_t;
subtype int956_t is signed(955 downto 0);
constant int956_t_SLV_LEN : integer := 956;
function int956_t_to_slv(x : int956_t) return std_logic_vector;
function slv_to_int956_t(x : std_logic_vector) return int956_t;
subtype uint957_t is unsigned(956 downto 0);
constant uint957_t_SLV_LEN : integer := 957;
function uint957_t_to_slv(x : uint957_t) return std_logic_vector;
function slv_to_uint957_t(x : std_logic_vector) return uint957_t;
subtype int957_t is signed(956 downto 0);
constant int957_t_SLV_LEN : integer := 957;
function int957_t_to_slv(x : int957_t) return std_logic_vector;
function slv_to_int957_t(x : std_logic_vector) return int957_t;
subtype uint958_t is unsigned(957 downto 0);
constant uint958_t_SLV_LEN : integer := 958;
function uint958_t_to_slv(x : uint958_t) return std_logic_vector;
function slv_to_uint958_t(x : std_logic_vector) return uint958_t;
subtype int958_t is signed(957 downto 0);
constant int958_t_SLV_LEN : integer := 958;
function int958_t_to_slv(x : int958_t) return std_logic_vector;
function slv_to_int958_t(x : std_logic_vector) return int958_t;
subtype uint959_t is unsigned(958 downto 0);
constant uint959_t_SLV_LEN : integer := 959;
function uint959_t_to_slv(x : uint959_t) return std_logic_vector;
function slv_to_uint959_t(x : std_logic_vector) return uint959_t;
subtype int959_t is signed(958 downto 0);
constant int959_t_SLV_LEN : integer := 959;
function int959_t_to_slv(x : int959_t) return std_logic_vector;
function slv_to_int959_t(x : std_logic_vector) return int959_t;
subtype uint960_t is unsigned(959 downto 0);
constant uint960_t_SLV_LEN : integer := 960;
function uint960_t_to_slv(x : uint960_t) return std_logic_vector;
function slv_to_uint960_t(x : std_logic_vector) return uint960_t;
subtype int960_t is signed(959 downto 0);
constant int960_t_SLV_LEN : integer := 960;
function int960_t_to_slv(x : int960_t) return std_logic_vector;
function slv_to_int960_t(x : std_logic_vector) return int960_t;
subtype uint961_t is unsigned(960 downto 0);
constant uint961_t_SLV_LEN : integer := 961;
function uint961_t_to_slv(x : uint961_t) return std_logic_vector;
function slv_to_uint961_t(x : std_logic_vector) return uint961_t;
subtype int961_t is signed(960 downto 0);
constant int961_t_SLV_LEN : integer := 961;
function int961_t_to_slv(x : int961_t) return std_logic_vector;
function slv_to_int961_t(x : std_logic_vector) return int961_t;
subtype uint962_t is unsigned(961 downto 0);
constant uint962_t_SLV_LEN : integer := 962;
function uint962_t_to_slv(x : uint962_t) return std_logic_vector;
function slv_to_uint962_t(x : std_logic_vector) return uint962_t;
subtype int962_t is signed(961 downto 0);
constant int962_t_SLV_LEN : integer := 962;
function int962_t_to_slv(x : int962_t) return std_logic_vector;
function slv_to_int962_t(x : std_logic_vector) return int962_t;
subtype uint963_t is unsigned(962 downto 0);
constant uint963_t_SLV_LEN : integer := 963;
function uint963_t_to_slv(x : uint963_t) return std_logic_vector;
function slv_to_uint963_t(x : std_logic_vector) return uint963_t;
subtype int963_t is signed(962 downto 0);
constant int963_t_SLV_LEN : integer := 963;
function int963_t_to_slv(x : int963_t) return std_logic_vector;
function slv_to_int963_t(x : std_logic_vector) return int963_t;
subtype uint964_t is unsigned(963 downto 0);
constant uint964_t_SLV_LEN : integer := 964;
function uint964_t_to_slv(x : uint964_t) return std_logic_vector;
function slv_to_uint964_t(x : std_logic_vector) return uint964_t;
subtype int964_t is signed(963 downto 0);
constant int964_t_SLV_LEN : integer := 964;
function int964_t_to_slv(x : int964_t) return std_logic_vector;
function slv_to_int964_t(x : std_logic_vector) return int964_t;
subtype uint965_t is unsigned(964 downto 0);
constant uint965_t_SLV_LEN : integer := 965;
function uint965_t_to_slv(x : uint965_t) return std_logic_vector;
function slv_to_uint965_t(x : std_logic_vector) return uint965_t;
subtype int965_t is signed(964 downto 0);
constant int965_t_SLV_LEN : integer := 965;
function int965_t_to_slv(x : int965_t) return std_logic_vector;
function slv_to_int965_t(x : std_logic_vector) return int965_t;
subtype uint966_t is unsigned(965 downto 0);
constant uint966_t_SLV_LEN : integer := 966;
function uint966_t_to_slv(x : uint966_t) return std_logic_vector;
function slv_to_uint966_t(x : std_logic_vector) return uint966_t;
subtype int966_t is signed(965 downto 0);
constant int966_t_SLV_LEN : integer := 966;
function int966_t_to_slv(x : int966_t) return std_logic_vector;
function slv_to_int966_t(x : std_logic_vector) return int966_t;
subtype uint967_t is unsigned(966 downto 0);
constant uint967_t_SLV_LEN : integer := 967;
function uint967_t_to_slv(x : uint967_t) return std_logic_vector;
function slv_to_uint967_t(x : std_logic_vector) return uint967_t;
subtype int967_t is signed(966 downto 0);
constant int967_t_SLV_LEN : integer := 967;
function int967_t_to_slv(x : int967_t) return std_logic_vector;
function slv_to_int967_t(x : std_logic_vector) return int967_t;
subtype uint968_t is unsigned(967 downto 0);
constant uint968_t_SLV_LEN : integer := 968;
function uint968_t_to_slv(x : uint968_t) return std_logic_vector;
function slv_to_uint968_t(x : std_logic_vector) return uint968_t;
subtype int968_t is signed(967 downto 0);
constant int968_t_SLV_LEN : integer := 968;
function int968_t_to_slv(x : int968_t) return std_logic_vector;
function slv_to_int968_t(x : std_logic_vector) return int968_t;
subtype uint969_t is unsigned(968 downto 0);
constant uint969_t_SLV_LEN : integer := 969;
function uint969_t_to_slv(x : uint969_t) return std_logic_vector;
function slv_to_uint969_t(x : std_logic_vector) return uint969_t;
subtype int969_t is signed(968 downto 0);
constant int969_t_SLV_LEN : integer := 969;
function int969_t_to_slv(x : int969_t) return std_logic_vector;
function slv_to_int969_t(x : std_logic_vector) return int969_t;
subtype uint970_t is unsigned(969 downto 0);
constant uint970_t_SLV_LEN : integer := 970;
function uint970_t_to_slv(x : uint970_t) return std_logic_vector;
function slv_to_uint970_t(x : std_logic_vector) return uint970_t;
subtype int970_t is signed(969 downto 0);
constant int970_t_SLV_LEN : integer := 970;
function int970_t_to_slv(x : int970_t) return std_logic_vector;
function slv_to_int970_t(x : std_logic_vector) return int970_t;
subtype uint971_t is unsigned(970 downto 0);
constant uint971_t_SLV_LEN : integer := 971;
function uint971_t_to_slv(x : uint971_t) return std_logic_vector;
function slv_to_uint971_t(x : std_logic_vector) return uint971_t;
subtype int971_t is signed(970 downto 0);
constant int971_t_SLV_LEN : integer := 971;
function int971_t_to_slv(x : int971_t) return std_logic_vector;
function slv_to_int971_t(x : std_logic_vector) return int971_t;
subtype uint972_t is unsigned(971 downto 0);
constant uint972_t_SLV_LEN : integer := 972;
function uint972_t_to_slv(x : uint972_t) return std_logic_vector;
function slv_to_uint972_t(x : std_logic_vector) return uint972_t;
subtype int972_t is signed(971 downto 0);
constant int972_t_SLV_LEN : integer := 972;
function int972_t_to_slv(x : int972_t) return std_logic_vector;
function slv_to_int972_t(x : std_logic_vector) return int972_t;
subtype uint973_t is unsigned(972 downto 0);
constant uint973_t_SLV_LEN : integer := 973;
function uint973_t_to_slv(x : uint973_t) return std_logic_vector;
function slv_to_uint973_t(x : std_logic_vector) return uint973_t;
subtype int973_t is signed(972 downto 0);
constant int973_t_SLV_LEN : integer := 973;
function int973_t_to_slv(x : int973_t) return std_logic_vector;
function slv_to_int973_t(x : std_logic_vector) return int973_t;
subtype uint974_t is unsigned(973 downto 0);
constant uint974_t_SLV_LEN : integer := 974;
function uint974_t_to_slv(x : uint974_t) return std_logic_vector;
function slv_to_uint974_t(x : std_logic_vector) return uint974_t;
subtype int974_t is signed(973 downto 0);
constant int974_t_SLV_LEN : integer := 974;
function int974_t_to_slv(x : int974_t) return std_logic_vector;
function slv_to_int974_t(x : std_logic_vector) return int974_t;
subtype uint975_t is unsigned(974 downto 0);
constant uint975_t_SLV_LEN : integer := 975;
function uint975_t_to_slv(x : uint975_t) return std_logic_vector;
function slv_to_uint975_t(x : std_logic_vector) return uint975_t;
subtype int975_t is signed(974 downto 0);
constant int975_t_SLV_LEN : integer := 975;
function int975_t_to_slv(x : int975_t) return std_logic_vector;
function slv_to_int975_t(x : std_logic_vector) return int975_t;
subtype uint976_t is unsigned(975 downto 0);
constant uint976_t_SLV_LEN : integer := 976;
function uint976_t_to_slv(x : uint976_t) return std_logic_vector;
function slv_to_uint976_t(x : std_logic_vector) return uint976_t;
subtype int976_t is signed(975 downto 0);
constant int976_t_SLV_LEN : integer := 976;
function int976_t_to_slv(x : int976_t) return std_logic_vector;
function slv_to_int976_t(x : std_logic_vector) return int976_t;
subtype uint977_t is unsigned(976 downto 0);
constant uint977_t_SLV_LEN : integer := 977;
function uint977_t_to_slv(x : uint977_t) return std_logic_vector;
function slv_to_uint977_t(x : std_logic_vector) return uint977_t;
subtype int977_t is signed(976 downto 0);
constant int977_t_SLV_LEN : integer := 977;
function int977_t_to_slv(x : int977_t) return std_logic_vector;
function slv_to_int977_t(x : std_logic_vector) return int977_t;
subtype uint978_t is unsigned(977 downto 0);
constant uint978_t_SLV_LEN : integer := 978;
function uint978_t_to_slv(x : uint978_t) return std_logic_vector;
function slv_to_uint978_t(x : std_logic_vector) return uint978_t;
subtype int978_t is signed(977 downto 0);
constant int978_t_SLV_LEN : integer := 978;
function int978_t_to_slv(x : int978_t) return std_logic_vector;
function slv_to_int978_t(x : std_logic_vector) return int978_t;
subtype uint979_t is unsigned(978 downto 0);
constant uint979_t_SLV_LEN : integer := 979;
function uint979_t_to_slv(x : uint979_t) return std_logic_vector;
function slv_to_uint979_t(x : std_logic_vector) return uint979_t;
subtype int979_t is signed(978 downto 0);
constant int979_t_SLV_LEN : integer := 979;
function int979_t_to_slv(x : int979_t) return std_logic_vector;
function slv_to_int979_t(x : std_logic_vector) return int979_t;
subtype uint980_t is unsigned(979 downto 0);
constant uint980_t_SLV_LEN : integer := 980;
function uint980_t_to_slv(x : uint980_t) return std_logic_vector;
function slv_to_uint980_t(x : std_logic_vector) return uint980_t;
subtype int980_t is signed(979 downto 0);
constant int980_t_SLV_LEN : integer := 980;
function int980_t_to_slv(x : int980_t) return std_logic_vector;
function slv_to_int980_t(x : std_logic_vector) return int980_t;
subtype uint981_t is unsigned(980 downto 0);
constant uint981_t_SLV_LEN : integer := 981;
function uint981_t_to_slv(x : uint981_t) return std_logic_vector;
function slv_to_uint981_t(x : std_logic_vector) return uint981_t;
subtype int981_t is signed(980 downto 0);
constant int981_t_SLV_LEN : integer := 981;
function int981_t_to_slv(x : int981_t) return std_logic_vector;
function slv_to_int981_t(x : std_logic_vector) return int981_t;
subtype uint982_t is unsigned(981 downto 0);
constant uint982_t_SLV_LEN : integer := 982;
function uint982_t_to_slv(x : uint982_t) return std_logic_vector;
function slv_to_uint982_t(x : std_logic_vector) return uint982_t;
subtype int982_t is signed(981 downto 0);
constant int982_t_SLV_LEN : integer := 982;
function int982_t_to_slv(x : int982_t) return std_logic_vector;
function slv_to_int982_t(x : std_logic_vector) return int982_t;
subtype uint983_t is unsigned(982 downto 0);
constant uint983_t_SLV_LEN : integer := 983;
function uint983_t_to_slv(x : uint983_t) return std_logic_vector;
function slv_to_uint983_t(x : std_logic_vector) return uint983_t;
subtype int983_t is signed(982 downto 0);
constant int983_t_SLV_LEN : integer := 983;
function int983_t_to_slv(x : int983_t) return std_logic_vector;
function slv_to_int983_t(x : std_logic_vector) return int983_t;
subtype uint984_t is unsigned(983 downto 0);
constant uint984_t_SLV_LEN : integer := 984;
function uint984_t_to_slv(x : uint984_t) return std_logic_vector;
function slv_to_uint984_t(x : std_logic_vector) return uint984_t;
subtype int984_t is signed(983 downto 0);
constant int984_t_SLV_LEN : integer := 984;
function int984_t_to_slv(x : int984_t) return std_logic_vector;
function slv_to_int984_t(x : std_logic_vector) return int984_t;
subtype uint985_t is unsigned(984 downto 0);
constant uint985_t_SLV_LEN : integer := 985;
function uint985_t_to_slv(x : uint985_t) return std_logic_vector;
function slv_to_uint985_t(x : std_logic_vector) return uint985_t;
subtype int985_t is signed(984 downto 0);
constant int985_t_SLV_LEN : integer := 985;
function int985_t_to_slv(x : int985_t) return std_logic_vector;
function slv_to_int985_t(x : std_logic_vector) return int985_t;
subtype uint986_t is unsigned(985 downto 0);
constant uint986_t_SLV_LEN : integer := 986;
function uint986_t_to_slv(x : uint986_t) return std_logic_vector;
function slv_to_uint986_t(x : std_logic_vector) return uint986_t;
subtype int986_t is signed(985 downto 0);
constant int986_t_SLV_LEN : integer := 986;
function int986_t_to_slv(x : int986_t) return std_logic_vector;
function slv_to_int986_t(x : std_logic_vector) return int986_t;
subtype uint987_t is unsigned(986 downto 0);
constant uint987_t_SLV_LEN : integer := 987;
function uint987_t_to_slv(x : uint987_t) return std_logic_vector;
function slv_to_uint987_t(x : std_logic_vector) return uint987_t;
subtype int987_t is signed(986 downto 0);
constant int987_t_SLV_LEN : integer := 987;
function int987_t_to_slv(x : int987_t) return std_logic_vector;
function slv_to_int987_t(x : std_logic_vector) return int987_t;
subtype uint988_t is unsigned(987 downto 0);
constant uint988_t_SLV_LEN : integer := 988;
function uint988_t_to_slv(x : uint988_t) return std_logic_vector;
function slv_to_uint988_t(x : std_logic_vector) return uint988_t;
subtype int988_t is signed(987 downto 0);
constant int988_t_SLV_LEN : integer := 988;
function int988_t_to_slv(x : int988_t) return std_logic_vector;
function slv_to_int988_t(x : std_logic_vector) return int988_t;
subtype uint989_t is unsigned(988 downto 0);
constant uint989_t_SLV_LEN : integer := 989;
function uint989_t_to_slv(x : uint989_t) return std_logic_vector;
function slv_to_uint989_t(x : std_logic_vector) return uint989_t;
subtype int989_t is signed(988 downto 0);
constant int989_t_SLV_LEN : integer := 989;
function int989_t_to_slv(x : int989_t) return std_logic_vector;
function slv_to_int989_t(x : std_logic_vector) return int989_t;
subtype uint990_t is unsigned(989 downto 0);
constant uint990_t_SLV_LEN : integer := 990;
function uint990_t_to_slv(x : uint990_t) return std_logic_vector;
function slv_to_uint990_t(x : std_logic_vector) return uint990_t;
subtype int990_t is signed(989 downto 0);
constant int990_t_SLV_LEN : integer := 990;
function int990_t_to_slv(x : int990_t) return std_logic_vector;
function slv_to_int990_t(x : std_logic_vector) return int990_t;
subtype uint991_t is unsigned(990 downto 0);
constant uint991_t_SLV_LEN : integer := 991;
function uint991_t_to_slv(x : uint991_t) return std_logic_vector;
function slv_to_uint991_t(x : std_logic_vector) return uint991_t;
subtype int991_t is signed(990 downto 0);
constant int991_t_SLV_LEN : integer := 991;
function int991_t_to_slv(x : int991_t) return std_logic_vector;
function slv_to_int991_t(x : std_logic_vector) return int991_t;
subtype uint992_t is unsigned(991 downto 0);
constant uint992_t_SLV_LEN : integer := 992;
function uint992_t_to_slv(x : uint992_t) return std_logic_vector;
function slv_to_uint992_t(x : std_logic_vector) return uint992_t;
subtype int992_t is signed(991 downto 0);
constant int992_t_SLV_LEN : integer := 992;
function int992_t_to_slv(x : int992_t) return std_logic_vector;
function slv_to_int992_t(x : std_logic_vector) return int992_t;
subtype uint993_t is unsigned(992 downto 0);
constant uint993_t_SLV_LEN : integer := 993;
function uint993_t_to_slv(x : uint993_t) return std_logic_vector;
function slv_to_uint993_t(x : std_logic_vector) return uint993_t;
subtype int993_t is signed(992 downto 0);
constant int993_t_SLV_LEN : integer := 993;
function int993_t_to_slv(x : int993_t) return std_logic_vector;
function slv_to_int993_t(x : std_logic_vector) return int993_t;
subtype uint994_t is unsigned(993 downto 0);
constant uint994_t_SLV_LEN : integer := 994;
function uint994_t_to_slv(x : uint994_t) return std_logic_vector;
function slv_to_uint994_t(x : std_logic_vector) return uint994_t;
subtype int994_t is signed(993 downto 0);
constant int994_t_SLV_LEN : integer := 994;
function int994_t_to_slv(x : int994_t) return std_logic_vector;
function slv_to_int994_t(x : std_logic_vector) return int994_t;
subtype uint995_t is unsigned(994 downto 0);
constant uint995_t_SLV_LEN : integer := 995;
function uint995_t_to_slv(x : uint995_t) return std_logic_vector;
function slv_to_uint995_t(x : std_logic_vector) return uint995_t;
subtype int995_t is signed(994 downto 0);
constant int995_t_SLV_LEN : integer := 995;
function int995_t_to_slv(x : int995_t) return std_logic_vector;
function slv_to_int995_t(x : std_logic_vector) return int995_t;
subtype uint996_t is unsigned(995 downto 0);
constant uint996_t_SLV_LEN : integer := 996;
function uint996_t_to_slv(x : uint996_t) return std_logic_vector;
function slv_to_uint996_t(x : std_logic_vector) return uint996_t;
subtype int996_t is signed(995 downto 0);
constant int996_t_SLV_LEN : integer := 996;
function int996_t_to_slv(x : int996_t) return std_logic_vector;
function slv_to_int996_t(x : std_logic_vector) return int996_t;
subtype uint997_t is unsigned(996 downto 0);
constant uint997_t_SLV_LEN : integer := 997;
function uint997_t_to_slv(x : uint997_t) return std_logic_vector;
function slv_to_uint997_t(x : std_logic_vector) return uint997_t;
subtype int997_t is signed(996 downto 0);
constant int997_t_SLV_LEN : integer := 997;
function int997_t_to_slv(x : int997_t) return std_logic_vector;
function slv_to_int997_t(x : std_logic_vector) return int997_t;
subtype uint998_t is unsigned(997 downto 0);
constant uint998_t_SLV_LEN : integer := 998;
function uint998_t_to_slv(x : uint998_t) return std_logic_vector;
function slv_to_uint998_t(x : std_logic_vector) return uint998_t;
subtype int998_t is signed(997 downto 0);
constant int998_t_SLV_LEN : integer := 998;
function int998_t_to_slv(x : int998_t) return std_logic_vector;
function slv_to_int998_t(x : std_logic_vector) return int998_t;
subtype uint999_t is unsigned(998 downto 0);
constant uint999_t_SLV_LEN : integer := 999;
function uint999_t_to_slv(x : uint999_t) return std_logic_vector;
function slv_to_uint999_t(x : std_logic_vector) return uint999_t;
subtype int999_t is signed(998 downto 0);
constant int999_t_SLV_LEN : integer := 999;
function int999_t_to_slv(x : int999_t) return std_logic_vector;
function slv_to_int999_t(x : std_logic_vector) return int999_t;
subtype uint1000_t is unsigned(999 downto 0);
constant uint1000_t_SLV_LEN : integer := 1000;
function uint1000_t_to_slv(x : uint1000_t) return std_logic_vector;
function slv_to_uint1000_t(x : std_logic_vector) return uint1000_t;
subtype int1000_t is signed(999 downto 0);
constant int1000_t_SLV_LEN : integer := 1000;
function int1000_t_to_slv(x : int1000_t) return std_logic_vector;
function slv_to_int1000_t(x : std_logic_vector) return int1000_t;
subtype uint1001_t is unsigned(1000 downto 0);
constant uint1001_t_SLV_LEN : integer := 1001;
function uint1001_t_to_slv(x : uint1001_t) return std_logic_vector;
function slv_to_uint1001_t(x : std_logic_vector) return uint1001_t;
subtype int1001_t is signed(1000 downto 0);
constant int1001_t_SLV_LEN : integer := 1001;
function int1001_t_to_slv(x : int1001_t) return std_logic_vector;
function slv_to_int1001_t(x : std_logic_vector) return int1001_t;
subtype uint1002_t is unsigned(1001 downto 0);
constant uint1002_t_SLV_LEN : integer := 1002;
function uint1002_t_to_slv(x : uint1002_t) return std_logic_vector;
function slv_to_uint1002_t(x : std_logic_vector) return uint1002_t;
subtype int1002_t is signed(1001 downto 0);
constant int1002_t_SLV_LEN : integer := 1002;
function int1002_t_to_slv(x : int1002_t) return std_logic_vector;
function slv_to_int1002_t(x : std_logic_vector) return int1002_t;
subtype uint1003_t is unsigned(1002 downto 0);
constant uint1003_t_SLV_LEN : integer := 1003;
function uint1003_t_to_slv(x : uint1003_t) return std_logic_vector;
function slv_to_uint1003_t(x : std_logic_vector) return uint1003_t;
subtype int1003_t is signed(1002 downto 0);
constant int1003_t_SLV_LEN : integer := 1003;
function int1003_t_to_slv(x : int1003_t) return std_logic_vector;
function slv_to_int1003_t(x : std_logic_vector) return int1003_t;
subtype uint1004_t is unsigned(1003 downto 0);
constant uint1004_t_SLV_LEN : integer := 1004;
function uint1004_t_to_slv(x : uint1004_t) return std_logic_vector;
function slv_to_uint1004_t(x : std_logic_vector) return uint1004_t;
subtype int1004_t is signed(1003 downto 0);
constant int1004_t_SLV_LEN : integer := 1004;
function int1004_t_to_slv(x : int1004_t) return std_logic_vector;
function slv_to_int1004_t(x : std_logic_vector) return int1004_t;
subtype uint1005_t is unsigned(1004 downto 0);
constant uint1005_t_SLV_LEN : integer := 1005;
function uint1005_t_to_slv(x : uint1005_t) return std_logic_vector;
function slv_to_uint1005_t(x : std_logic_vector) return uint1005_t;
subtype int1005_t is signed(1004 downto 0);
constant int1005_t_SLV_LEN : integer := 1005;
function int1005_t_to_slv(x : int1005_t) return std_logic_vector;
function slv_to_int1005_t(x : std_logic_vector) return int1005_t;
subtype uint1006_t is unsigned(1005 downto 0);
constant uint1006_t_SLV_LEN : integer := 1006;
function uint1006_t_to_slv(x : uint1006_t) return std_logic_vector;
function slv_to_uint1006_t(x : std_logic_vector) return uint1006_t;
subtype int1006_t is signed(1005 downto 0);
constant int1006_t_SLV_LEN : integer := 1006;
function int1006_t_to_slv(x : int1006_t) return std_logic_vector;
function slv_to_int1006_t(x : std_logic_vector) return int1006_t;
subtype uint1007_t is unsigned(1006 downto 0);
constant uint1007_t_SLV_LEN : integer := 1007;
function uint1007_t_to_slv(x : uint1007_t) return std_logic_vector;
function slv_to_uint1007_t(x : std_logic_vector) return uint1007_t;
subtype int1007_t is signed(1006 downto 0);
constant int1007_t_SLV_LEN : integer := 1007;
function int1007_t_to_slv(x : int1007_t) return std_logic_vector;
function slv_to_int1007_t(x : std_logic_vector) return int1007_t;
subtype uint1008_t is unsigned(1007 downto 0);
constant uint1008_t_SLV_LEN : integer := 1008;
function uint1008_t_to_slv(x : uint1008_t) return std_logic_vector;
function slv_to_uint1008_t(x : std_logic_vector) return uint1008_t;
subtype int1008_t is signed(1007 downto 0);
constant int1008_t_SLV_LEN : integer := 1008;
function int1008_t_to_slv(x : int1008_t) return std_logic_vector;
function slv_to_int1008_t(x : std_logic_vector) return int1008_t;
subtype uint1009_t is unsigned(1008 downto 0);
constant uint1009_t_SLV_LEN : integer := 1009;
function uint1009_t_to_slv(x : uint1009_t) return std_logic_vector;
function slv_to_uint1009_t(x : std_logic_vector) return uint1009_t;
subtype int1009_t is signed(1008 downto 0);
constant int1009_t_SLV_LEN : integer := 1009;
function int1009_t_to_slv(x : int1009_t) return std_logic_vector;
function slv_to_int1009_t(x : std_logic_vector) return int1009_t;
subtype uint1010_t is unsigned(1009 downto 0);
constant uint1010_t_SLV_LEN : integer := 1010;
function uint1010_t_to_slv(x : uint1010_t) return std_logic_vector;
function slv_to_uint1010_t(x : std_logic_vector) return uint1010_t;
subtype int1010_t is signed(1009 downto 0);
constant int1010_t_SLV_LEN : integer := 1010;
function int1010_t_to_slv(x : int1010_t) return std_logic_vector;
function slv_to_int1010_t(x : std_logic_vector) return int1010_t;
subtype uint1011_t is unsigned(1010 downto 0);
constant uint1011_t_SLV_LEN : integer := 1011;
function uint1011_t_to_slv(x : uint1011_t) return std_logic_vector;
function slv_to_uint1011_t(x : std_logic_vector) return uint1011_t;
subtype int1011_t is signed(1010 downto 0);
constant int1011_t_SLV_LEN : integer := 1011;
function int1011_t_to_slv(x : int1011_t) return std_logic_vector;
function slv_to_int1011_t(x : std_logic_vector) return int1011_t;
subtype uint1012_t is unsigned(1011 downto 0);
constant uint1012_t_SLV_LEN : integer := 1012;
function uint1012_t_to_slv(x : uint1012_t) return std_logic_vector;
function slv_to_uint1012_t(x : std_logic_vector) return uint1012_t;
subtype int1012_t is signed(1011 downto 0);
constant int1012_t_SLV_LEN : integer := 1012;
function int1012_t_to_slv(x : int1012_t) return std_logic_vector;
function slv_to_int1012_t(x : std_logic_vector) return int1012_t;
subtype uint1013_t is unsigned(1012 downto 0);
constant uint1013_t_SLV_LEN : integer := 1013;
function uint1013_t_to_slv(x : uint1013_t) return std_logic_vector;
function slv_to_uint1013_t(x : std_logic_vector) return uint1013_t;
subtype int1013_t is signed(1012 downto 0);
constant int1013_t_SLV_LEN : integer := 1013;
function int1013_t_to_slv(x : int1013_t) return std_logic_vector;
function slv_to_int1013_t(x : std_logic_vector) return int1013_t;
subtype uint1014_t is unsigned(1013 downto 0);
constant uint1014_t_SLV_LEN : integer := 1014;
function uint1014_t_to_slv(x : uint1014_t) return std_logic_vector;
function slv_to_uint1014_t(x : std_logic_vector) return uint1014_t;
subtype int1014_t is signed(1013 downto 0);
constant int1014_t_SLV_LEN : integer := 1014;
function int1014_t_to_slv(x : int1014_t) return std_logic_vector;
function slv_to_int1014_t(x : std_logic_vector) return int1014_t;
subtype uint1015_t is unsigned(1014 downto 0);
constant uint1015_t_SLV_LEN : integer := 1015;
function uint1015_t_to_slv(x : uint1015_t) return std_logic_vector;
function slv_to_uint1015_t(x : std_logic_vector) return uint1015_t;
subtype int1015_t is signed(1014 downto 0);
constant int1015_t_SLV_LEN : integer := 1015;
function int1015_t_to_slv(x : int1015_t) return std_logic_vector;
function slv_to_int1015_t(x : std_logic_vector) return int1015_t;
subtype uint1016_t is unsigned(1015 downto 0);
constant uint1016_t_SLV_LEN : integer := 1016;
function uint1016_t_to_slv(x : uint1016_t) return std_logic_vector;
function slv_to_uint1016_t(x : std_logic_vector) return uint1016_t;
subtype int1016_t is signed(1015 downto 0);
constant int1016_t_SLV_LEN : integer := 1016;
function int1016_t_to_slv(x : int1016_t) return std_logic_vector;
function slv_to_int1016_t(x : std_logic_vector) return int1016_t;
subtype uint1017_t is unsigned(1016 downto 0);
constant uint1017_t_SLV_LEN : integer := 1017;
function uint1017_t_to_slv(x : uint1017_t) return std_logic_vector;
function slv_to_uint1017_t(x : std_logic_vector) return uint1017_t;
subtype int1017_t is signed(1016 downto 0);
constant int1017_t_SLV_LEN : integer := 1017;
function int1017_t_to_slv(x : int1017_t) return std_logic_vector;
function slv_to_int1017_t(x : std_logic_vector) return int1017_t;
subtype uint1018_t is unsigned(1017 downto 0);
constant uint1018_t_SLV_LEN : integer := 1018;
function uint1018_t_to_slv(x : uint1018_t) return std_logic_vector;
function slv_to_uint1018_t(x : std_logic_vector) return uint1018_t;
subtype int1018_t is signed(1017 downto 0);
constant int1018_t_SLV_LEN : integer := 1018;
function int1018_t_to_slv(x : int1018_t) return std_logic_vector;
function slv_to_int1018_t(x : std_logic_vector) return int1018_t;
subtype uint1019_t is unsigned(1018 downto 0);
constant uint1019_t_SLV_LEN : integer := 1019;
function uint1019_t_to_slv(x : uint1019_t) return std_logic_vector;
function slv_to_uint1019_t(x : std_logic_vector) return uint1019_t;
subtype int1019_t is signed(1018 downto 0);
constant int1019_t_SLV_LEN : integer := 1019;
function int1019_t_to_slv(x : int1019_t) return std_logic_vector;
function slv_to_int1019_t(x : std_logic_vector) return int1019_t;
subtype uint1020_t is unsigned(1019 downto 0);
constant uint1020_t_SLV_LEN : integer := 1020;
function uint1020_t_to_slv(x : uint1020_t) return std_logic_vector;
function slv_to_uint1020_t(x : std_logic_vector) return uint1020_t;
subtype int1020_t is signed(1019 downto 0);
constant int1020_t_SLV_LEN : integer := 1020;
function int1020_t_to_slv(x : int1020_t) return std_logic_vector;
function slv_to_int1020_t(x : std_logic_vector) return int1020_t;
subtype uint1021_t is unsigned(1020 downto 0);
constant uint1021_t_SLV_LEN : integer := 1021;
function uint1021_t_to_slv(x : uint1021_t) return std_logic_vector;
function slv_to_uint1021_t(x : std_logic_vector) return uint1021_t;
subtype int1021_t is signed(1020 downto 0);
constant int1021_t_SLV_LEN : integer := 1021;
function int1021_t_to_slv(x : int1021_t) return std_logic_vector;
function slv_to_int1021_t(x : std_logic_vector) return int1021_t;
subtype uint1022_t is unsigned(1021 downto 0);
constant uint1022_t_SLV_LEN : integer := 1022;
function uint1022_t_to_slv(x : uint1022_t) return std_logic_vector;
function slv_to_uint1022_t(x : std_logic_vector) return uint1022_t;
subtype int1022_t is signed(1021 downto 0);
constant int1022_t_SLV_LEN : integer := 1022;
function int1022_t_to_slv(x : int1022_t) return std_logic_vector;
function slv_to_int1022_t(x : std_logic_vector) return int1022_t;
subtype uint1023_t is unsigned(1022 downto 0);
constant uint1023_t_SLV_LEN : integer := 1023;
function uint1023_t_to_slv(x : uint1023_t) return std_logic_vector;
function slv_to_uint1023_t(x : std_logic_vector) return uint1023_t;
subtype int1023_t is signed(1022 downto 0);
constant int1023_t_SLV_LEN : integer := 1023;
function int1023_t_to_slv(x : int1023_t) return std_logic_vector;
function slv_to_int1023_t(x : std_logic_vector) return int1023_t;
subtype uint1024_t is unsigned(1023 downto 0);
constant uint1024_t_SLV_LEN : integer := 1024;
function uint1024_t_to_slv(x : uint1024_t) return std_logic_vector;
function slv_to_uint1024_t(x : std_logic_vector) return uint1024_t;
subtype int1024_t is signed(1023 downto 0);
constant int1024_t_SLV_LEN : integer := 1024;
function int1024_t_to_slv(x : int1024_t) return std_logic_vector;
function slv_to_int1024_t(x : std_logic_vector) return int1024_t;
subtype uint1025_t is unsigned(1024 downto 0);
constant uint1025_t_SLV_LEN : integer := 1025;
function uint1025_t_to_slv(x : uint1025_t) return std_logic_vector;
function slv_to_uint1025_t(x : std_logic_vector) return uint1025_t;
subtype int1025_t is signed(1024 downto 0);
constant int1025_t_SLV_LEN : integer := 1025;
function int1025_t_to_slv(x : int1025_t) return std_logic_vector;
function slv_to_int1025_t(x : std_logic_vector) return int1025_t;
subtype uint1026_t is unsigned(1025 downto 0);
constant uint1026_t_SLV_LEN : integer := 1026;
function uint1026_t_to_slv(x : uint1026_t) return std_logic_vector;
function slv_to_uint1026_t(x : std_logic_vector) return uint1026_t;
subtype int1026_t is signed(1025 downto 0);
constant int1026_t_SLV_LEN : integer := 1026;
function int1026_t_to_slv(x : int1026_t) return std_logic_vector;
function slv_to_int1026_t(x : std_logic_vector) return int1026_t;
subtype uint1027_t is unsigned(1026 downto 0);
constant uint1027_t_SLV_LEN : integer := 1027;
function uint1027_t_to_slv(x : uint1027_t) return std_logic_vector;
function slv_to_uint1027_t(x : std_logic_vector) return uint1027_t;
subtype int1027_t is signed(1026 downto 0);
constant int1027_t_SLV_LEN : integer := 1027;
function int1027_t_to_slv(x : int1027_t) return std_logic_vector;
function slv_to_int1027_t(x : std_logic_vector) return int1027_t;
subtype uint1028_t is unsigned(1027 downto 0);
constant uint1028_t_SLV_LEN : integer := 1028;
function uint1028_t_to_slv(x : uint1028_t) return std_logic_vector;
function slv_to_uint1028_t(x : std_logic_vector) return uint1028_t;
subtype int1028_t is signed(1027 downto 0);
constant int1028_t_SLV_LEN : integer := 1028;
function int1028_t_to_slv(x : int1028_t) return std_logic_vector;
function slv_to_int1028_t(x : std_logic_vector) return int1028_t;
subtype uint1029_t is unsigned(1028 downto 0);
constant uint1029_t_SLV_LEN : integer := 1029;
function uint1029_t_to_slv(x : uint1029_t) return std_logic_vector;
function slv_to_uint1029_t(x : std_logic_vector) return uint1029_t;
subtype int1029_t is signed(1028 downto 0);
constant int1029_t_SLV_LEN : integer := 1029;
function int1029_t_to_slv(x : int1029_t) return std_logic_vector;
function slv_to_int1029_t(x : std_logic_vector) return int1029_t;
subtype uint1030_t is unsigned(1029 downto 0);
constant uint1030_t_SLV_LEN : integer := 1030;
function uint1030_t_to_slv(x : uint1030_t) return std_logic_vector;
function slv_to_uint1030_t(x : std_logic_vector) return uint1030_t;
subtype int1030_t is signed(1029 downto 0);
constant int1030_t_SLV_LEN : integer := 1030;
function int1030_t_to_slv(x : int1030_t) return std_logic_vector;
function slv_to_int1030_t(x : std_logic_vector) return int1030_t;
subtype uint1031_t is unsigned(1030 downto 0);
constant uint1031_t_SLV_LEN : integer := 1031;
function uint1031_t_to_slv(x : uint1031_t) return std_logic_vector;
function slv_to_uint1031_t(x : std_logic_vector) return uint1031_t;
subtype int1031_t is signed(1030 downto 0);
constant int1031_t_SLV_LEN : integer := 1031;
function int1031_t_to_slv(x : int1031_t) return std_logic_vector;
function slv_to_int1031_t(x : std_logic_vector) return int1031_t;
subtype uint1032_t is unsigned(1031 downto 0);
constant uint1032_t_SLV_LEN : integer := 1032;
function uint1032_t_to_slv(x : uint1032_t) return std_logic_vector;
function slv_to_uint1032_t(x : std_logic_vector) return uint1032_t;
subtype int1032_t is signed(1031 downto 0);
constant int1032_t_SLV_LEN : integer := 1032;
function int1032_t_to_slv(x : int1032_t) return std_logic_vector;
function slv_to_int1032_t(x : std_logic_vector) return int1032_t;
subtype uint1033_t is unsigned(1032 downto 0);
constant uint1033_t_SLV_LEN : integer := 1033;
function uint1033_t_to_slv(x : uint1033_t) return std_logic_vector;
function slv_to_uint1033_t(x : std_logic_vector) return uint1033_t;
subtype int1033_t is signed(1032 downto 0);
constant int1033_t_SLV_LEN : integer := 1033;
function int1033_t_to_slv(x : int1033_t) return std_logic_vector;
function slv_to_int1033_t(x : std_logic_vector) return int1033_t;
subtype uint1034_t is unsigned(1033 downto 0);
constant uint1034_t_SLV_LEN : integer := 1034;
function uint1034_t_to_slv(x : uint1034_t) return std_logic_vector;
function slv_to_uint1034_t(x : std_logic_vector) return uint1034_t;
subtype int1034_t is signed(1033 downto 0);
constant int1034_t_SLV_LEN : integer := 1034;
function int1034_t_to_slv(x : int1034_t) return std_logic_vector;
function slv_to_int1034_t(x : std_logic_vector) return int1034_t;
subtype uint1035_t is unsigned(1034 downto 0);
constant uint1035_t_SLV_LEN : integer := 1035;
function uint1035_t_to_slv(x : uint1035_t) return std_logic_vector;
function slv_to_uint1035_t(x : std_logic_vector) return uint1035_t;
subtype int1035_t is signed(1034 downto 0);
constant int1035_t_SLV_LEN : integer := 1035;
function int1035_t_to_slv(x : int1035_t) return std_logic_vector;
function slv_to_int1035_t(x : std_logic_vector) return int1035_t;
subtype uint1036_t is unsigned(1035 downto 0);
constant uint1036_t_SLV_LEN : integer := 1036;
function uint1036_t_to_slv(x : uint1036_t) return std_logic_vector;
function slv_to_uint1036_t(x : std_logic_vector) return uint1036_t;
subtype int1036_t is signed(1035 downto 0);
constant int1036_t_SLV_LEN : integer := 1036;
function int1036_t_to_slv(x : int1036_t) return std_logic_vector;
function slv_to_int1036_t(x : std_logic_vector) return int1036_t;
subtype uint1037_t is unsigned(1036 downto 0);
constant uint1037_t_SLV_LEN : integer := 1037;
function uint1037_t_to_slv(x : uint1037_t) return std_logic_vector;
function slv_to_uint1037_t(x : std_logic_vector) return uint1037_t;
subtype int1037_t is signed(1036 downto 0);
constant int1037_t_SLV_LEN : integer := 1037;
function int1037_t_to_slv(x : int1037_t) return std_logic_vector;
function slv_to_int1037_t(x : std_logic_vector) return int1037_t;
subtype uint1038_t is unsigned(1037 downto 0);
constant uint1038_t_SLV_LEN : integer := 1038;
function uint1038_t_to_slv(x : uint1038_t) return std_logic_vector;
function slv_to_uint1038_t(x : std_logic_vector) return uint1038_t;
subtype int1038_t is signed(1037 downto 0);
constant int1038_t_SLV_LEN : integer := 1038;
function int1038_t_to_slv(x : int1038_t) return std_logic_vector;
function slv_to_int1038_t(x : std_logic_vector) return int1038_t;
subtype uint1039_t is unsigned(1038 downto 0);
constant uint1039_t_SLV_LEN : integer := 1039;
function uint1039_t_to_slv(x : uint1039_t) return std_logic_vector;
function slv_to_uint1039_t(x : std_logic_vector) return uint1039_t;
subtype int1039_t is signed(1038 downto 0);
constant int1039_t_SLV_LEN : integer := 1039;
function int1039_t_to_slv(x : int1039_t) return std_logic_vector;
function slv_to_int1039_t(x : std_logic_vector) return int1039_t;
subtype uint1040_t is unsigned(1039 downto 0);
constant uint1040_t_SLV_LEN : integer := 1040;
function uint1040_t_to_slv(x : uint1040_t) return std_logic_vector;
function slv_to_uint1040_t(x : std_logic_vector) return uint1040_t;
subtype int1040_t is signed(1039 downto 0);
constant int1040_t_SLV_LEN : integer := 1040;
function int1040_t_to_slv(x : int1040_t) return std_logic_vector;
function slv_to_int1040_t(x : std_logic_vector) return int1040_t;
subtype uint1041_t is unsigned(1040 downto 0);
constant uint1041_t_SLV_LEN : integer := 1041;
function uint1041_t_to_slv(x : uint1041_t) return std_logic_vector;
function slv_to_uint1041_t(x : std_logic_vector) return uint1041_t;
subtype int1041_t is signed(1040 downto 0);
constant int1041_t_SLV_LEN : integer := 1041;
function int1041_t_to_slv(x : int1041_t) return std_logic_vector;
function slv_to_int1041_t(x : std_logic_vector) return int1041_t;
subtype uint1042_t is unsigned(1041 downto 0);
constant uint1042_t_SLV_LEN : integer := 1042;
function uint1042_t_to_slv(x : uint1042_t) return std_logic_vector;
function slv_to_uint1042_t(x : std_logic_vector) return uint1042_t;
subtype int1042_t is signed(1041 downto 0);
constant int1042_t_SLV_LEN : integer := 1042;
function int1042_t_to_slv(x : int1042_t) return std_logic_vector;
function slv_to_int1042_t(x : std_logic_vector) return int1042_t;
subtype uint1043_t is unsigned(1042 downto 0);
constant uint1043_t_SLV_LEN : integer := 1043;
function uint1043_t_to_slv(x : uint1043_t) return std_logic_vector;
function slv_to_uint1043_t(x : std_logic_vector) return uint1043_t;
subtype int1043_t is signed(1042 downto 0);
constant int1043_t_SLV_LEN : integer := 1043;
function int1043_t_to_slv(x : int1043_t) return std_logic_vector;
function slv_to_int1043_t(x : std_logic_vector) return int1043_t;
subtype uint1044_t is unsigned(1043 downto 0);
constant uint1044_t_SLV_LEN : integer := 1044;
function uint1044_t_to_slv(x : uint1044_t) return std_logic_vector;
function slv_to_uint1044_t(x : std_logic_vector) return uint1044_t;
subtype int1044_t is signed(1043 downto 0);
constant int1044_t_SLV_LEN : integer := 1044;
function int1044_t_to_slv(x : int1044_t) return std_logic_vector;
function slv_to_int1044_t(x : std_logic_vector) return int1044_t;
subtype uint1045_t is unsigned(1044 downto 0);
constant uint1045_t_SLV_LEN : integer := 1045;
function uint1045_t_to_slv(x : uint1045_t) return std_logic_vector;
function slv_to_uint1045_t(x : std_logic_vector) return uint1045_t;
subtype int1045_t is signed(1044 downto 0);
constant int1045_t_SLV_LEN : integer := 1045;
function int1045_t_to_slv(x : int1045_t) return std_logic_vector;
function slv_to_int1045_t(x : std_logic_vector) return int1045_t;
subtype uint1046_t is unsigned(1045 downto 0);
constant uint1046_t_SLV_LEN : integer := 1046;
function uint1046_t_to_slv(x : uint1046_t) return std_logic_vector;
function slv_to_uint1046_t(x : std_logic_vector) return uint1046_t;
subtype int1046_t is signed(1045 downto 0);
constant int1046_t_SLV_LEN : integer := 1046;
function int1046_t_to_slv(x : int1046_t) return std_logic_vector;
function slv_to_int1046_t(x : std_logic_vector) return int1046_t;
subtype uint1047_t is unsigned(1046 downto 0);
constant uint1047_t_SLV_LEN : integer := 1047;
function uint1047_t_to_slv(x : uint1047_t) return std_logic_vector;
function slv_to_uint1047_t(x : std_logic_vector) return uint1047_t;
subtype int1047_t is signed(1046 downto 0);
constant int1047_t_SLV_LEN : integer := 1047;
function int1047_t_to_slv(x : int1047_t) return std_logic_vector;
function slv_to_int1047_t(x : std_logic_vector) return int1047_t;
subtype uint1048_t is unsigned(1047 downto 0);
constant uint1048_t_SLV_LEN : integer := 1048;
function uint1048_t_to_slv(x : uint1048_t) return std_logic_vector;
function slv_to_uint1048_t(x : std_logic_vector) return uint1048_t;
subtype int1048_t is signed(1047 downto 0);
constant int1048_t_SLV_LEN : integer := 1048;
function int1048_t_to_slv(x : int1048_t) return std_logic_vector;
function slv_to_int1048_t(x : std_logic_vector) return int1048_t;
subtype uint1049_t is unsigned(1048 downto 0);
constant uint1049_t_SLV_LEN : integer := 1049;
function uint1049_t_to_slv(x : uint1049_t) return std_logic_vector;
function slv_to_uint1049_t(x : std_logic_vector) return uint1049_t;
subtype int1049_t is signed(1048 downto 0);
constant int1049_t_SLV_LEN : integer := 1049;
function int1049_t_to_slv(x : int1049_t) return std_logic_vector;
function slv_to_int1049_t(x : std_logic_vector) return int1049_t;
subtype uint1050_t is unsigned(1049 downto 0);
constant uint1050_t_SLV_LEN : integer := 1050;
function uint1050_t_to_slv(x : uint1050_t) return std_logic_vector;
function slv_to_uint1050_t(x : std_logic_vector) return uint1050_t;
subtype int1050_t is signed(1049 downto 0);
constant int1050_t_SLV_LEN : integer := 1050;
function int1050_t_to_slv(x : int1050_t) return std_logic_vector;
function slv_to_int1050_t(x : std_logic_vector) return int1050_t;
subtype uint1051_t is unsigned(1050 downto 0);
constant uint1051_t_SLV_LEN : integer := 1051;
function uint1051_t_to_slv(x : uint1051_t) return std_logic_vector;
function slv_to_uint1051_t(x : std_logic_vector) return uint1051_t;
subtype int1051_t is signed(1050 downto 0);
constant int1051_t_SLV_LEN : integer := 1051;
function int1051_t_to_slv(x : int1051_t) return std_logic_vector;
function slv_to_int1051_t(x : std_logic_vector) return int1051_t;
subtype uint1052_t is unsigned(1051 downto 0);
constant uint1052_t_SLV_LEN : integer := 1052;
function uint1052_t_to_slv(x : uint1052_t) return std_logic_vector;
function slv_to_uint1052_t(x : std_logic_vector) return uint1052_t;
subtype int1052_t is signed(1051 downto 0);
constant int1052_t_SLV_LEN : integer := 1052;
function int1052_t_to_slv(x : int1052_t) return std_logic_vector;
function slv_to_int1052_t(x : std_logic_vector) return int1052_t;
subtype uint1053_t is unsigned(1052 downto 0);
constant uint1053_t_SLV_LEN : integer := 1053;
function uint1053_t_to_slv(x : uint1053_t) return std_logic_vector;
function slv_to_uint1053_t(x : std_logic_vector) return uint1053_t;
subtype int1053_t is signed(1052 downto 0);
constant int1053_t_SLV_LEN : integer := 1053;
function int1053_t_to_slv(x : int1053_t) return std_logic_vector;
function slv_to_int1053_t(x : std_logic_vector) return int1053_t;
subtype uint1054_t is unsigned(1053 downto 0);
constant uint1054_t_SLV_LEN : integer := 1054;
function uint1054_t_to_slv(x : uint1054_t) return std_logic_vector;
function slv_to_uint1054_t(x : std_logic_vector) return uint1054_t;
subtype int1054_t is signed(1053 downto 0);
constant int1054_t_SLV_LEN : integer := 1054;
function int1054_t_to_slv(x : int1054_t) return std_logic_vector;
function slv_to_int1054_t(x : std_logic_vector) return int1054_t;
subtype uint1055_t is unsigned(1054 downto 0);
constant uint1055_t_SLV_LEN : integer := 1055;
function uint1055_t_to_slv(x : uint1055_t) return std_logic_vector;
function slv_to_uint1055_t(x : std_logic_vector) return uint1055_t;
subtype int1055_t is signed(1054 downto 0);
constant int1055_t_SLV_LEN : integer := 1055;
function int1055_t_to_slv(x : int1055_t) return std_logic_vector;
function slv_to_int1055_t(x : std_logic_vector) return int1055_t;
subtype uint1056_t is unsigned(1055 downto 0);
constant uint1056_t_SLV_LEN : integer := 1056;
function uint1056_t_to_slv(x : uint1056_t) return std_logic_vector;
function slv_to_uint1056_t(x : std_logic_vector) return uint1056_t;
subtype int1056_t is signed(1055 downto 0);
constant int1056_t_SLV_LEN : integer := 1056;
function int1056_t_to_slv(x : int1056_t) return std_logic_vector;
function slv_to_int1056_t(x : std_logic_vector) return int1056_t;
subtype uint1057_t is unsigned(1056 downto 0);
constant uint1057_t_SLV_LEN : integer := 1057;
function uint1057_t_to_slv(x : uint1057_t) return std_logic_vector;
function slv_to_uint1057_t(x : std_logic_vector) return uint1057_t;
subtype int1057_t is signed(1056 downto 0);
constant int1057_t_SLV_LEN : integer := 1057;
function int1057_t_to_slv(x : int1057_t) return std_logic_vector;
function slv_to_int1057_t(x : std_logic_vector) return int1057_t;
subtype uint1058_t is unsigned(1057 downto 0);
constant uint1058_t_SLV_LEN : integer := 1058;
function uint1058_t_to_slv(x : uint1058_t) return std_logic_vector;
function slv_to_uint1058_t(x : std_logic_vector) return uint1058_t;
subtype int1058_t is signed(1057 downto 0);
constant int1058_t_SLV_LEN : integer := 1058;
function int1058_t_to_slv(x : int1058_t) return std_logic_vector;
function slv_to_int1058_t(x : std_logic_vector) return int1058_t;
subtype uint1059_t is unsigned(1058 downto 0);
constant uint1059_t_SLV_LEN : integer := 1059;
function uint1059_t_to_slv(x : uint1059_t) return std_logic_vector;
function slv_to_uint1059_t(x : std_logic_vector) return uint1059_t;
subtype int1059_t is signed(1058 downto 0);
constant int1059_t_SLV_LEN : integer := 1059;
function int1059_t_to_slv(x : int1059_t) return std_logic_vector;
function slv_to_int1059_t(x : std_logic_vector) return int1059_t;
subtype uint1060_t is unsigned(1059 downto 0);
constant uint1060_t_SLV_LEN : integer := 1060;
function uint1060_t_to_slv(x : uint1060_t) return std_logic_vector;
function slv_to_uint1060_t(x : std_logic_vector) return uint1060_t;
subtype int1060_t is signed(1059 downto 0);
constant int1060_t_SLV_LEN : integer := 1060;
function int1060_t_to_slv(x : int1060_t) return std_logic_vector;
function slv_to_int1060_t(x : std_logic_vector) return int1060_t;
subtype uint1061_t is unsigned(1060 downto 0);
constant uint1061_t_SLV_LEN : integer := 1061;
function uint1061_t_to_slv(x : uint1061_t) return std_logic_vector;
function slv_to_uint1061_t(x : std_logic_vector) return uint1061_t;
subtype int1061_t is signed(1060 downto 0);
constant int1061_t_SLV_LEN : integer := 1061;
function int1061_t_to_slv(x : int1061_t) return std_logic_vector;
function slv_to_int1061_t(x : std_logic_vector) return int1061_t;
subtype uint1062_t is unsigned(1061 downto 0);
constant uint1062_t_SLV_LEN : integer := 1062;
function uint1062_t_to_slv(x : uint1062_t) return std_logic_vector;
function slv_to_uint1062_t(x : std_logic_vector) return uint1062_t;
subtype int1062_t is signed(1061 downto 0);
constant int1062_t_SLV_LEN : integer := 1062;
function int1062_t_to_slv(x : int1062_t) return std_logic_vector;
function slv_to_int1062_t(x : std_logic_vector) return int1062_t;
subtype uint1063_t is unsigned(1062 downto 0);
constant uint1063_t_SLV_LEN : integer := 1063;
function uint1063_t_to_slv(x : uint1063_t) return std_logic_vector;
function slv_to_uint1063_t(x : std_logic_vector) return uint1063_t;
subtype int1063_t is signed(1062 downto 0);
constant int1063_t_SLV_LEN : integer := 1063;
function int1063_t_to_slv(x : int1063_t) return std_logic_vector;
function slv_to_int1063_t(x : std_logic_vector) return int1063_t;
subtype uint1064_t is unsigned(1063 downto 0);
constant uint1064_t_SLV_LEN : integer := 1064;
function uint1064_t_to_slv(x : uint1064_t) return std_logic_vector;
function slv_to_uint1064_t(x : std_logic_vector) return uint1064_t;
subtype int1064_t is signed(1063 downto 0);
constant int1064_t_SLV_LEN : integer := 1064;
function int1064_t_to_slv(x : int1064_t) return std_logic_vector;
function slv_to_int1064_t(x : std_logic_vector) return int1064_t;
subtype uint1065_t is unsigned(1064 downto 0);
constant uint1065_t_SLV_LEN : integer := 1065;
function uint1065_t_to_slv(x : uint1065_t) return std_logic_vector;
function slv_to_uint1065_t(x : std_logic_vector) return uint1065_t;
subtype int1065_t is signed(1064 downto 0);
constant int1065_t_SLV_LEN : integer := 1065;
function int1065_t_to_slv(x : int1065_t) return std_logic_vector;
function slv_to_int1065_t(x : std_logic_vector) return int1065_t;
subtype uint1066_t is unsigned(1065 downto 0);
constant uint1066_t_SLV_LEN : integer := 1066;
function uint1066_t_to_slv(x : uint1066_t) return std_logic_vector;
function slv_to_uint1066_t(x : std_logic_vector) return uint1066_t;
subtype int1066_t is signed(1065 downto 0);
constant int1066_t_SLV_LEN : integer := 1066;
function int1066_t_to_slv(x : int1066_t) return std_logic_vector;
function slv_to_int1066_t(x : std_logic_vector) return int1066_t;
subtype uint1067_t is unsigned(1066 downto 0);
constant uint1067_t_SLV_LEN : integer := 1067;
function uint1067_t_to_slv(x : uint1067_t) return std_logic_vector;
function slv_to_uint1067_t(x : std_logic_vector) return uint1067_t;
subtype int1067_t is signed(1066 downto 0);
constant int1067_t_SLV_LEN : integer := 1067;
function int1067_t_to_slv(x : int1067_t) return std_logic_vector;
function slv_to_int1067_t(x : std_logic_vector) return int1067_t;
subtype uint1068_t is unsigned(1067 downto 0);
constant uint1068_t_SLV_LEN : integer := 1068;
function uint1068_t_to_slv(x : uint1068_t) return std_logic_vector;
function slv_to_uint1068_t(x : std_logic_vector) return uint1068_t;
subtype int1068_t is signed(1067 downto 0);
constant int1068_t_SLV_LEN : integer := 1068;
function int1068_t_to_slv(x : int1068_t) return std_logic_vector;
function slv_to_int1068_t(x : std_logic_vector) return int1068_t;
subtype uint1069_t is unsigned(1068 downto 0);
constant uint1069_t_SLV_LEN : integer := 1069;
function uint1069_t_to_slv(x : uint1069_t) return std_logic_vector;
function slv_to_uint1069_t(x : std_logic_vector) return uint1069_t;
subtype int1069_t is signed(1068 downto 0);
constant int1069_t_SLV_LEN : integer := 1069;
function int1069_t_to_slv(x : int1069_t) return std_logic_vector;
function slv_to_int1069_t(x : std_logic_vector) return int1069_t;
subtype uint1070_t is unsigned(1069 downto 0);
constant uint1070_t_SLV_LEN : integer := 1070;
function uint1070_t_to_slv(x : uint1070_t) return std_logic_vector;
function slv_to_uint1070_t(x : std_logic_vector) return uint1070_t;
subtype int1070_t is signed(1069 downto 0);
constant int1070_t_SLV_LEN : integer := 1070;
function int1070_t_to_slv(x : int1070_t) return std_logic_vector;
function slv_to_int1070_t(x : std_logic_vector) return int1070_t;
subtype uint1071_t is unsigned(1070 downto 0);
constant uint1071_t_SLV_LEN : integer := 1071;
function uint1071_t_to_slv(x : uint1071_t) return std_logic_vector;
function slv_to_uint1071_t(x : std_logic_vector) return uint1071_t;
subtype int1071_t is signed(1070 downto 0);
constant int1071_t_SLV_LEN : integer := 1071;
function int1071_t_to_slv(x : int1071_t) return std_logic_vector;
function slv_to_int1071_t(x : std_logic_vector) return int1071_t;
subtype uint1072_t is unsigned(1071 downto 0);
constant uint1072_t_SLV_LEN : integer := 1072;
function uint1072_t_to_slv(x : uint1072_t) return std_logic_vector;
function slv_to_uint1072_t(x : std_logic_vector) return uint1072_t;
subtype int1072_t is signed(1071 downto 0);
constant int1072_t_SLV_LEN : integer := 1072;
function int1072_t_to_slv(x : int1072_t) return std_logic_vector;
function slv_to_int1072_t(x : std_logic_vector) return int1072_t;
subtype uint1073_t is unsigned(1072 downto 0);
constant uint1073_t_SLV_LEN : integer := 1073;
function uint1073_t_to_slv(x : uint1073_t) return std_logic_vector;
function slv_to_uint1073_t(x : std_logic_vector) return uint1073_t;
subtype int1073_t is signed(1072 downto 0);
constant int1073_t_SLV_LEN : integer := 1073;
function int1073_t_to_slv(x : int1073_t) return std_logic_vector;
function slv_to_int1073_t(x : std_logic_vector) return int1073_t;
subtype uint1074_t is unsigned(1073 downto 0);
constant uint1074_t_SLV_LEN : integer := 1074;
function uint1074_t_to_slv(x : uint1074_t) return std_logic_vector;
function slv_to_uint1074_t(x : std_logic_vector) return uint1074_t;
subtype int1074_t is signed(1073 downto 0);
constant int1074_t_SLV_LEN : integer := 1074;
function int1074_t_to_slv(x : int1074_t) return std_logic_vector;
function slv_to_int1074_t(x : std_logic_vector) return int1074_t;
subtype uint1075_t is unsigned(1074 downto 0);
constant uint1075_t_SLV_LEN : integer := 1075;
function uint1075_t_to_slv(x : uint1075_t) return std_logic_vector;
function slv_to_uint1075_t(x : std_logic_vector) return uint1075_t;
subtype int1075_t is signed(1074 downto 0);
constant int1075_t_SLV_LEN : integer := 1075;
function int1075_t_to_slv(x : int1075_t) return std_logic_vector;
function slv_to_int1075_t(x : std_logic_vector) return int1075_t;
subtype uint1076_t is unsigned(1075 downto 0);
constant uint1076_t_SLV_LEN : integer := 1076;
function uint1076_t_to_slv(x : uint1076_t) return std_logic_vector;
function slv_to_uint1076_t(x : std_logic_vector) return uint1076_t;
subtype int1076_t is signed(1075 downto 0);
constant int1076_t_SLV_LEN : integer := 1076;
function int1076_t_to_slv(x : int1076_t) return std_logic_vector;
function slv_to_int1076_t(x : std_logic_vector) return int1076_t;
subtype uint1077_t is unsigned(1076 downto 0);
constant uint1077_t_SLV_LEN : integer := 1077;
function uint1077_t_to_slv(x : uint1077_t) return std_logic_vector;
function slv_to_uint1077_t(x : std_logic_vector) return uint1077_t;
subtype int1077_t is signed(1076 downto 0);
constant int1077_t_SLV_LEN : integer := 1077;
function int1077_t_to_slv(x : int1077_t) return std_logic_vector;
function slv_to_int1077_t(x : std_logic_vector) return int1077_t;
subtype uint1078_t is unsigned(1077 downto 0);
constant uint1078_t_SLV_LEN : integer := 1078;
function uint1078_t_to_slv(x : uint1078_t) return std_logic_vector;
function slv_to_uint1078_t(x : std_logic_vector) return uint1078_t;
subtype int1078_t is signed(1077 downto 0);
constant int1078_t_SLV_LEN : integer := 1078;
function int1078_t_to_slv(x : int1078_t) return std_logic_vector;
function slv_to_int1078_t(x : std_logic_vector) return int1078_t;
subtype uint1079_t is unsigned(1078 downto 0);
constant uint1079_t_SLV_LEN : integer := 1079;
function uint1079_t_to_slv(x : uint1079_t) return std_logic_vector;
function slv_to_uint1079_t(x : std_logic_vector) return uint1079_t;
subtype int1079_t is signed(1078 downto 0);
constant int1079_t_SLV_LEN : integer := 1079;
function int1079_t_to_slv(x : int1079_t) return std_logic_vector;
function slv_to_int1079_t(x : std_logic_vector) return int1079_t;
subtype uint1080_t is unsigned(1079 downto 0);
constant uint1080_t_SLV_LEN : integer := 1080;
function uint1080_t_to_slv(x : uint1080_t) return std_logic_vector;
function slv_to_uint1080_t(x : std_logic_vector) return uint1080_t;
subtype int1080_t is signed(1079 downto 0);
constant int1080_t_SLV_LEN : integer := 1080;
function int1080_t_to_slv(x : int1080_t) return std_logic_vector;
function slv_to_int1080_t(x : std_logic_vector) return int1080_t;
subtype uint1081_t is unsigned(1080 downto 0);
constant uint1081_t_SLV_LEN : integer := 1081;
function uint1081_t_to_slv(x : uint1081_t) return std_logic_vector;
function slv_to_uint1081_t(x : std_logic_vector) return uint1081_t;
subtype int1081_t is signed(1080 downto 0);
constant int1081_t_SLV_LEN : integer := 1081;
function int1081_t_to_slv(x : int1081_t) return std_logic_vector;
function slv_to_int1081_t(x : std_logic_vector) return int1081_t;
subtype uint1082_t is unsigned(1081 downto 0);
constant uint1082_t_SLV_LEN : integer := 1082;
function uint1082_t_to_slv(x : uint1082_t) return std_logic_vector;
function slv_to_uint1082_t(x : std_logic_vector) return uint1082_t;
subtype int1082_t is signed(1081 downto 0);
constant int1082_t_SLV_LEN : integer := 1082;
function int1082_t_to_slv(x : int1082_t) return std_logic_vector;
function slv_to_int1082_t(x : std_logic_vector) return int1082_t;
subtype uint1083_t is unsigned(1082 downto 0);
constant uint1083_t_SLV_LEN : integer := 1083;
function uint1083_t_to_slv(x : uint1083_t) return std_logic_vector;
function slv_to_uint1083_t(x : std_logic_vector) return uint1083_t;
subtype int1083_t is signed(1082 downto 0);
constant int1083_t_SLV_LEN : integer := 1083;
function int1083_t_to_slv(x : int1083_t) return std_logic_vector;
function slv_to_int1083_t(x : std_logic_vector) return int1083_t;
subtype uint1084_t is unsigned(1083 downto 0);
constant uint1084_t_SLV_LEN : integer := 1084;
function uint1084_t_to_slv(x : uint1084_t) return std_logic_vector;
function slv_to_uint1084_t(x : std_logic_vector) return uint1084_t;
subtype int1084_t is signed(1083 downto 0);
constant int1084_t_SLV_LEN : integer := 1084;
function int1084_t_to_slv(x : int1084_t) return std_logic_vector;
function slv_to_int1084_t(x : std_logic_vector) return int1084_t;
subtype uint1085_t is unsigned(1084 downto 0);
constant uint1085_t_SLV_LEN : integer := 1085;
function uint1085_t_to_slv(x : uint1085_t) return std_logic_vector;
function slv_to_uint1085_t(x : std_logic_vector) return uint1085_t;
subtype int1085_t is signed(1084 downto 0);
constant int1085_t_SLV_LEN : integer := 1085;
function int1085_t_to_slv(x : int1085_t) return std_logic_vector;
function slv_to_int1085_t(x : std_logic_vector) return int1085_t;
subtype uint1086_t is unsigned(1085 downto 0);
constant uint1086_t_SLV_LEN : integer := 1086;
function uint1086_t_to_slv(x : uint1086_t) return std_logic_vector;
function slv_to_uint1086_t(x : std_logic_vector) return uint1086_t;
subtype int1086_t is signed(1085 downto 0);
constant int1086_t_SLV_LEN : integer := 1086;
function int1086_t_to_slv(x : int1086_t) return std_logic_vector;
function slv_to_int1086_t(x : std_logic_vector) return int1086_t;
subtype uint1087_t is unsigned(1086 downto 0);
constant uint1087_t_SLV_LEN : integer := 1087;
function uint1087_t_to_slv(x : uint1087_t) return std_logic_vector;
function slv_to_uint1087_t(x : std_logic_vector) return uint1087_t;
subtype int1087_t is signed(1086 downto 0);
constant int1087_t_SLV_LEN : integer := 1087;
function int1087_t_to_slv(x : int1087_t) return std_logic_vector;
function slv_to_int1087_t(x : std_logic_vector) return int1087_t;
subtype uint1088_t is unsigned(1087 downto 0);
constant uint1088_t_SLV_LEN : integer := 1088;
function uint1088_t_to_slv(x : uint1088_t) return std_logic_vector;
function slv_to_uint1088_t(x : std_logic_vector) return uint1088_t;
subtype int1088_t is signed(1087 downto 0);
constant int1088_t_SLV_LEN : integer := 1088;
function int1088_t_to_slv(x : int1088_t) return std_logic_vector;
function slv_to_int1088_t(x : std_logic_vector) return int1088_t;
subtype uint1089_t is unsigned(1088 downto 0);
constant uint1089_t_SLV_LEN : integer := 1089;
function uint1089_t_to_slv(x : uint1089_t) return std_logic_vector;
function slv_to_uint1089_t(x : std_logic_vector) return uint1089_t;
subtype int1089_t is signed(1088 downto 0);
constant int1089_t_SLV_LEN : integer := 1089;
function int1089_t_to_slv(x : int1089_t) return std_logic_vector;
function slv_to_int1089_t(x : std_logic_vector) return int1089_t;
subtype uint1090_t is unsigned(1089 downto 0);
constant uint1090_t_SLV_LEN : integer := 1090;
function uint1090_t_to_slv(x : uint1090_t) return std_logic_vector;
function slv_to_uint1090_t(x : std_logic_vector) return uint1090_t;
subtype int1090_t is signed(1089 downto 0);
constant int1090_t_SLV_LEN : integer := 1090;
function int1090_t_to_slv(x : int1090_t) return std_logic_vector;
function slv_to_int1090_t(x : std_logic_vector) return int1090_t;
subtype uint1091_t is unsigned(1090 downto 0);
constant uint1091_t_SLV_LEN : integer := 1091;
function uint1091_t_to_slv(x : uint1091_t) return std_logic_vector;
function slv_to_uint1091_t(x : std_logic_vector) return uint1091_t;
subtype int1091_t is signed(1090 downto 0);
constant int1091_t_SLV_LEN : integer := 1091;
function int1091_t_to_slv(x : int1091_t) return std_logic_vector;
function slv_to_int1091_t(x : std_logic_vector) return int1091_t;
subtype uint1092_t is unsigned(1091 downto 0);
constant uint1092_t_SLV_LEN : integer := 1092;
function uint1092_t_to_slv(x : uint1092_t) return std_logic_vector;
function slv_to_uint1092_t(x : std_logic_vector) return uint1092_t;
subtype int1092_t is signed(1091 downto 0);
constant int1092_t_SLV_LEN : integer := 1092;
function int1092_t_to_slv(x : int1092_t) return std_logic_vector;
function slv_to_int1092_t(x : std_logic_vector) return int1092_t;
subtype uint1093_t is unsigned(1092 downto 0);
constant uint1093_t_SLV_LEN : integer := 1093;
function uint1093_t_to_slv(x : uint1093_t) return std_logic_vector;
function slv_to_uint1093_t(x : std_logic_vector) return uint1093_t;
subtype int1093_t is signed(1092 downto 0);
constant int1093_t_SLV_LEN : integer := 1093;
function int1093_t_to_slv(x : int1093_t) return std_logic_vector;
function slv_to_int1093_t(x : std_logic_vector) return int1093_t;
subtype uint1094_t is unsigned(1093 downto 0);
constant uint1094_t_SLV_LEN : integer := 1094;
function uint1094_t_to_slv(x : uint1094_t) return std_logic_vector;
function slv_to_uint1094_t(x : std_logic_vector) return uint1094_t;
subtype int1094_t is signed(1093 downto 0);
constant int1094_t_SLV_LEN : integer := 1094;
function int1094_t_to_slv(x : int1094_t) return std_logic_vector;
function slv_to_int1094_t(x : std_logic_vector) return int1094_t;
subtype uint1095_t is unsigned(1094 downto 0);
constant uint1095_t_SLV_LEN : integer := 1095;
function uint1095_t_to_slv(x : uint1095_t) return std_logic_vector;
function slv_to_uint1095_t(x : std_logic_vector) return uint1095_t;
subtype int1095_t is signed(1094 downto 0);
constant int1095_t_SLV_LEN : integer := 1095;
function int1095_t_to_slv(x : int1095_t) return std_logic_vector;
function slv_to_int1095_t(x : std_logic_vector) return int1095_t;
subtype uint1096_t is unsigned(1095 downto 0);
constant uint1096_t_SLV_LEN : integer := 1096;
function uint1096_t_to_slv(x : uint1096_t) return std_logic_vector;
function slv_to_uint1096_t(x : std_logic_vector) return uint1096_t;
subtype int1096_t is signed(1095 downto 0);
constant int1096_t_SLV_LEN : integer := 1096;
function int1096_t_to_slv(x : int1096_t) return std_logic_vector;
function slv_to_int1096_t(x : std_logic_vector) return int1096_t;
subtype uint1097_t is unsigned(1096 downto 0);
constant uint1097_t_SLV_LEN : integer := 1097;
function uint1097_t_to_slv(x : uint1097_t) return std_logic_vector;
function slv_to_uint1097_t(x : std_logic_vector) return uint1097_t;
subtype int1097_t is signed(1096 downto 0);
constant int1097_t_SLV_LEN : integer := 1097;
function int1097_t_to_slv(x : int1097_t) return std_logic_vector;
function slv_to_int1097_t(x : std_logic_vector) return int1097_t;
subtype uint1098_t is unsigned(1097 downto 0);
constant uint1098_t_SLV_LEN : integer := 1098;
function uint1098_t_to_slv(x : uint1098_t) return std_logic_vector;
function slv_to_uint1098_t(x : std_logic_vector) return uint1098_t;
subtype int1098_t is signed(1097 downto 0);
constant int1098_t_SLV_LEN : integer := 1098;
function int1098_t_to_slv(x : int1098_t) return std_logic_vector;
function slv_to_int1098_t(x : std_logic_vector) return int1098_t;
subtype uint1099_t is unsigned(1098 downto 0);
constant uint1099_t_SLV_LEN : integer := 1099;
function uint1099_t_to_slv(x : uint1099_t) return std_logic_vector;
function slv_to_uint1099_t(x : std_logic_vector) return uint1099_t;
subtype int1099_t is signed(1098 downto 0);
constant int1099_t_SLV_LEN : integer := 1099;
function int1099_t_to_slv(x : int1099_t) return std_logic_vector;
function slv_to_int1099_t(x : std_logic_vector) return int1099_t;
subtype uint1100_t is unsigned(1099 downto 0);
constant uint1100_t_SLV_LEN : integer := 1100;
function uint1100_t_to_slv(x : uint1100_t) return std_logic_vector;
function slv_to_uint1100_t(x : std_logic_vector) return uint1100_t;
subtype int1100_t is signed(1099 downto 0);
constant int1100_t_SLV_LEN : integer := 1100;
function int1100_t_to_slv(x : int1100_t) return std_logic_vector;
function slv_to_int1100_t(x : std_logic_vector) return int1100_t;
subtype uint1101_t is unsigned(1100 downto 0);
constant uint1101_t_SLV_LEN : integer := 1101;
function uint1101_t_to_slv(x : uint1101_t) return std_logic_vector;
function slv_to_uint1101_t(x : std_logic_vector) return uint1101_t;
subtype int1101_t is signed(1100 downto 0);
constant int1101_t_SLV_LEN : integer := 1101;
function int1101_t_to_slv(x : int1101_t) return std_logic_vector;
function slv_to_int1101_t(x : std_logic_vector) return int1101_t;
subtype uint1102_t is unsigned(1101 downto 0);
constant uint1102_t_SLV_LEN : integer := 1102;
function uint1102_t_to_slv(x : uint1102_t) return std_logic_vector;
function slv_to_uint1102_t(x : std_logic_vector) return uint1102_t;
subtype int1102_t is signed(1101 downto 0);
constant int1102_t_SLV_LEN : integer := 1102;
function int1102_t_to_slv(x : int1102_t) return std_logic_vector;
function slv_to_int1102_t(x : std_logic_vector) return int1102_t;
subtype uint1103_t is unsigned(1102 downto 0);
constant uint1103_t_SLV_LEN : integer := 1103;
function uint1103_t_to_slv(x : uint1103_t) return std_logic_vector;
function slv_to_uint1103_t(x : std_logic_vector) return uint1103_t;
subtype int1103_t is signed(1102 downto 0);
constant int1103_t_SLV_LEN : integer := 1103;
function int1103_t_to_slv(x : int1103_t) return std_logic_vector;
function slv_to_int1103_t(x : std_logic_vector) return int1103_t;
subtype uint1104_t is unsigned(1103 downto 0);
constant uint1104_t_SLV_LEN : integer := 1104;
function uint1104_t_to_slv(x : uint1104_t) return std_logic_vector;
function slv_to_uint1104_t(x : std_logic_vector) return uint1104_t;
subtype int1104_t is signed(1103 downto 0);
constant int1104_t_SLV_LEN : integer := 1104;
function int1104_t_to_slv(x : int1104_t) return std_logic_vector;
function slv_to_int1104_t(x : std_logic_vector) return int1104_t;
subtype uint1105_t is unsigned(1104 downto 0);
constant uint1105_t_SLV_LEN : integer := 1105;
function uint1105_t_to_slv(x : uint1105_t) return std_logic_vector;
function slv_to_uint1105_t(x : std_logic_vector) return uint1105_t;
subtype int1105_t is signed(1104 downto 0);
constant int1105_t_SLV_LEN : integer := 1105;
function int1105_t_to_slv(x : int1105_t) return std_logic_vector;
function slv_to_int1105_t(x : std_logic_vector) return int1105_t;
subtype uint1106_t is unsigned(1105 downto 0);
constant uint1106_t_SLV_LEN : integer := 1106;
function uint1106_t_to_slv(x : uint1106_t) return std_logic_vector;
function slv_to_uint1106_t(x : std_logic_vector) return uint1106_t;
subtype int1106_t is signed(1105 downto 0);
constant int1106_t_SLV_LEN : integer := 1106;
function int1106_t_to_slv(x : int1106_t) return std_logic_vector;
function slv_to_int1106_t(x : std_logic_vector) return int1106_t;
subtype uint1107_t is unsigned(1106 downto 0);
constant uint1107_t_SLV_LEN : integer := 1107;
function uint1107_t_to_slv(x : uint1107_t) return std_logic_vector;
function slv_to_uint1107_t(x : std_logic_vector) return uint1107_t;
subtype int1107_t is signed(1106 downto 0);
constant int1107_t_SLV_LEN : integer := 1107;
function int1107_t_to_slv(x : int1107_t) return std_logic_vector;
function slv_to_int1107_t(x : std_logic_vector) return int1107_t;
subtype uint1108_t is unsigned(1107 downto 0);
constant uint1108_t_SLV_LEN : integer := 1108;
function uint1108_t_to_slv(x : uint1108_t) return std_logic_vector;
function slv_to_uint1108_t(x : std_logic_vector) return uint1108_t;
subtype int1108_t is signed(1107 downto 0);
constant int1108_t_SLV_LEN : integer := 1108;
function int1108_t_to_slv(x : int1108_t) return std_logic_vector;
function slv_to_int1108_t(x : std_logic_vector) return int1108_t;
subtype uint1109_t is unsigned(1108 downto 0);
constant uint1109_t_SLV_LEN : integer := 1109;
function uint1109_t_to_slv(x : uint1109_t) return std_logic_vector;
function slv_to_uint1109_t(x : std_logic_vector) return uint1109_t;
subtype int1109_t is signed(1108 downto 0);
constant int1109_t_SLV_LEN : integer := 1109;
function int1109_t_to_slv(x : int1109_t) return std_logic_vector;
function slv_to_int1109_t(x : std_logic_vector) return int1109_t;
subtype uint1110_t is unsigned(1109 downto 0);
constant uint1110_t_SLV_LEN : integer := 1110;
function uint1110_t_to_slv(x : uint1110_t) return std_logic_vector;
function slv_to_uint1110_t(x : std_logic_vector) return uint1110_t;
subtype int1110_t is signed(1109 downto 0);
constant int1110_t_SLV_LEN : integer := 1110;
function int1110_t_to_slv(x : int1110_t) return std_logic_vector;
function slv_to_int1110_t(x : std_logic_vector) return int1110_t;
subtype uint1111_t is unsigned(1110 downto 0);
constant uint1111_t_SLV_LEN : integer := 1111;
function uint1111_t_to_slv(x : uint1111_t) return std_logic_vector;
function slv_to_uint1111_t(x : std_logic_vector) return uint1111_t;
subtype int1111_t is signed(1110 downto 0);
constant int1111_t_SLV_LEN : integer := 1111;
function int1111_t_to_slv(x : int1111_t) return std_logic_vector;
function slv_to_int1111_t(x : std_logic_vector) return int1111_t;
subtype uint1112_t is unsigned(1111 downto 0);
constant uint1112_t_SLV_LEN : integer := 1112;
function uint1112_t_to_slv(x : uint1112_t) return std_logic_vector;
function slv_to_uint1112_t(x : std_logic_vector) return uint1112_t;
subtype int1112_t is signed(1111 downto 0);
constant int1112_t_SLV_LEN : integer := 1112;
function int1112_t_to_slv(x : int1112_t) return std_logic_vector;
function slv_to_int1112_t(x : std_logic_vector) return int1112_t;
subtype uint1113_t is unsigned(1112 downto 0);
constant uint1113_t_SLV_LEN : integer := 1113;
function uint1113_t_to_slv(x : uint1113_t) return std_logic_vector;
function slv_to_uint1113_t(x : std_logic_vector) return uint1113_t;
subtype int1113_t is signed(1112 downto 0);
constant int1113_t_SLV_LEN : integer := 1113;
function int1113_t_to_slv(x : int1113_t) return std_logic_vector;
function slv_to_int1113_t(x : std_logic_vector) return int1113_t;
subtype uint1114_t is unsigned(1113 downto 0);
constant uint1114_t_SLV_LEN : integer := 1114;
function uint1114_t_to_slv(x : uint1114_t) return std_logic_vector;
function slv_to_uint1114_t(x : std_logic_vector) return uint1114_t;
subtype int1114_t is signed(1113 downto 0);
constant int1114_t_SLV_LEN : integer := 1114;
function int1114_t_to_slv(x : int1114_t) return std_logic_vector;
function slv_to_int1114_t(x : std_logic_vector) return int1114_t;
subtype uint1115_t is unsigned(1114 downto 0);
constant uint1115_t_SLV_LEN : integer := 1115;
function uint1115_t_to_slv(x : uint1115_t) return std_logic_vector;
function slv_to_uint1115_t(x : std_logic_vector) return uint1115_t;
subtype int1115_t is signed(1114 downto 0);
constant int1115_t_SLV_LEN : integer := 1115;
function int1115_t_to_slv(x : int1115_t) return std_logic_vector;
function slv_to_int1115_t(x : std_logic_vector) return int1115_t;
subtype uint1116_t is unsigned(1115 downto 0);
constant uint1116_t_SLV_LEN : integer := 1116;
function uint1116_t_to_slv(x : uint1116_t) return std_logic_vector;
function slv_to_uint1116_t(x : std_logic_vector) return uint1116_t;
subtype int1116_t is signed(1115 downto 0);
constant int1116_t_SLV_LEN : integer := 1116;
function int1116_t_to_slv(x : int1116_t) return std_logic_vector;
function slv_to_int1116_t(x : std_logic_vector) return int1116_t;
subtype uint1117_t is unsigned(1116 downto 0);
constant uint1117_t_SLV_LEN : integer := 1117;
function uint1117_t_to_slv(x : uint1117_t) return std_logic_vector;
function slv_to_uint1117_t(x : std_logic_vector) return uint1117_t;
subtype int1117_t is signed(1116 downto 0);
constant int1117_t_SLV_LEN : integer := 1117;
function int1117_t_to_slv(x : int1117_t) return std_logic_vector;
function slv_to_int1117_t(x : std_logic_vector) return int1117_t;
subtype uint1118_t is unsigned(1117 downto 0);
constant uint1118_t_SLV_LEN : integer := 1118;
function uint1118_t_to_slv(x : uint1118_t) return std_logic_vector;
function slv_to_uint1118_t(x : std_logic_vector) return uint1118_t;
subtype int1118_t is signed(1117 downto 0);
constant int1118_t_SLV_LEN : integer := 1118;
function int1118_t_to_slv(x : int1118_t) return std_logic_vector;
function slv_to_int1118_t(x : std_logic_vector) return int1118_t;
subtype uint1119_t is unsigned(1118 downto 0);
constant uint1119_t_SLV_LEN : integer := 1119;
function uint1119_t_to_slv(x : uint1119_t) return std_logic_vector;
function slv_to_uint1119_t(x : std_logic_vector) return uint1119_t;
subtype int1119_t is signed(1118 downto 0);
constant int1119_t_SLV_LEN : integer := 1119;
function int1119_t_to_slv(x : int1119_t) return std_logic_vector;
function slv_to_int1119_t(x : std_logic_vector) return int1119_t;
subtype uint1120_t is unsigned(1119 downto 0);
constant uint1120_t_SLV_LEN : integer := 1120;
function uint1120_t_to_slv(x : uint1120_t) return std_logic_vector;
function slv_to_uint1120_t(x : std_logic_vector) return uint1120_t;
subtype int1120_t is signed(1119 downto 0);
constant int1120_t_SLV_LEN : integer := 1120;
function int1120_t_to_slv(x : int1120_t) return std_logic_vector;
function slv_to_int1120_t(x : std_logic_vector) return int1120_t;
subtype uint1121_t is unsigned(1120 downto 0);
constant uint1121_t_SLV_LEN : integer := 1121;
function uint1121_t_to_slv(x : uint1121_t) return std_logic_vector;
function slv_to_uint1121_t(x : std_logic_vector) return uint1121_t;
subtype int1121_t is signed(1120 downto 0);
constant int1121_t_SLV_LEN : integer := 1121;
function int1121_t_to_slv(x : int1121_t) return std_logic_vector;
function slv_to_int1121_t(x : std_logic_vector) return int1121_t;
subtype uint1122_t is unsigned(1121 downto 0);
constant uint1122_t_SLV_LEN : integer := 1122;
function uint1122_t_to_slv(x : uint1122_t) return std_logic_vector;
function slv_to_uint1122_t(x : std_logic_vector) return uint1122_t;
subtype int1122_t is signed(1121 downto 0);
constant int1122_t_SLV_LEN : integer := 1122;
function int1122_t_to_slv(x : int1122_t) return std_logic_vector;
function slv_to_int1122_t(x : std_logic_vector) return int1122_t;
subtype uint1123_t is unsigned(1122 downto 0);
constant uint1123_t_SLV_LEN : integer := 1123;
function uint1123_t_to_slv(x : uint1123_t) return std_logic_vector;
function slv_to_uint1123_t(x : std_logic_vector) return uint1123_t;
subtype int1123_t is signed(1122 downto 0);
constant int1123_t_SLV_LEN : integer := 1123;
function int1123_t_to_slv(x : int1123_t) return std_logic_vector;
function slv_to_int1123_t(x : std_logic_vector) return int1123_t;
subtype uint1124_t is unsigned(1123 downto 0);
constant uint1124_t_SLV_LEN : integer := 1124;
function uint1124_t_to_slv(x : uint1124_t) return std_logic_vector;
function slv_to_uint1124_t(x : std_logic_vector) return uint1124_t;
subtype int1124_t is signed(1123 downto 0);
constant int1124_t_SLV_LEN : integer := 1124;
function int1124_t_to_slv(x : int1124_t) return std_logic_vector;
function slv_to_int1124_t(x : std_logic_vector) return int1124_t;
subtype uint1125_t is unsigned(1124 downto 0);
constant uint1125_t_SLV_LEN : integer := 1125;
function uint1125_t_to_slv(x : uint1125_t) return std_logic_vector;
function slv_to_uint1125_t(x : std_logic_vector) return uint1125_t;
subtype int1125_t is signed(1124 downto 0);
constant int1125_t_SLV_LEN : integer := 1125;
function int1125_t_to_slv(x : int1125_t) return std_logic_vector;
function slv_to_int1125_t(x : std_logic_vector) return int1125_t;
subtype uint1126_t is unsigned(1125 downto 0);
constant uint1126_t_SLV_LEN : integer := 1126;
function uint1126_t_to_slv(x : uint1126_t) return std_logic_vector;
function slv_to_uint1126_t(x : std_logic_vector) return uint1126_t;
subtype int1126_t is signed(1125 downto 0);
constant int1126_t_SLV_LEN : integer := 1126;
function int1126_t_to_slv(x : int1126_t) return std_logic_vector;
function slv_to_int1126_t(x : std_logic_vector) return int1126_t;
subtype uint1127_t is unsigned(1126 downto 0);
constant uint1127_t_SLV_LEN : integer := 1127;
function uint1127_t_to_slv(x : uint1127_t) return std_logic_vector;
function slv_to_uint1127_t(x : std_logic_vector) return uint1127_t;
subtype int1127_t is signed(1126 downto 0);
constant int1127_t_SLV_LEN : integer := 1127;
function int1127_t_to_slv(x : int1127_t) return std_logic_vector;
function slv_to_int1127_t(x : std_logic_vector) return int1127_t;
subtype uint1128_t is unsigned(1127 downto 0);
constant uint1128_t_SLV_LEN : integer := 1128;
function uint1128_t_to_slv(x : uint1128_t) return std_logic_vector;
function slv_to_uint1128_t(x : std_logic_vector) return uint1128_t;
subtype int1128_t is signed(1127 downto 0);
constant int1128_t_SLV_LEN : integer := 1128;
function int1128_t_to_slv(x : int1128_t) return std_logic_vector;
function slv_to_int1128_t(x : std_logic_vector) return int1128_t;
subtype uint1129_t is unsigned(1128 downto 0);
constant uint1129_t_SLV_LEN : integer := 1129;
function uint1129_t_to_slv(x : uint1129_t) return std_logic_vector;
function slv_to_uint1129_t(x : std_logic_vector) return uint1129_t;
subtype int1129_t is signed(1128 downto 0);
constant int1129_t_SLV_LEN : integer := 1129;
function int1129_t_to_slv(x : int1129_t) return std_logic_vector;
function slv_to_int1129_t(x : std_logic_vector) return int1129_t;
subtype uint1130_t is unsigned(1129 downto 0);
constant uint1130_t_SLV_LEN : integer := 1130;
function uint1130_t_to_slv(x : uint1130_t) return std_logic_vector;
function slv_to_uint1130_t(x : std_logic_vector) return uint1130_t;
subtype int1130_t is signed(1129 downto 0);
constant int1130_t_SLV_LEN : integer := 1130;
function int1130_t_to_slv(x : int1130_t) return std_logic_vector;
function slv_to_int1130_t(x : std_logic_vector) return int1130_t;
subtype uint1131_t is unsigned(1130 downto 0);
constant uint1131_t_SLV_LEN : integer := 1131;
function uint1131_t_to_slv(x : uint1131_t) return std_logic_vector;
function slv_to_uint1131_t(x : std_logic_vector) return uint1131_t;
subtype int1131_t is signed(1130 downto 0);
constant int1131_t_SLV_LEN : integer := 1131;
function int1131_t_to_slv(x : int1131_t) return std_logic_vector;
function slv_to_int1131_t(x : std_logic_vector) return int1131_t;
subtype uint1132_t is unsigned(1131 downto 0);
constant uint1132_t_SLV_LEN : integer := 1132;
function uint1132_t_to_slv(x : uint1132_t) return std_logic_vector;
function slv_to_uint1132_t(x : std_logic_vector) return uint1132_t;
subtype int1132_t is signed(1131 downto 0);
constant int1132_t_SLV_LEN : integer := 1132;
function int1132_t_to_slv(x : int1132_t) return std_logic_vector;
function slv_to_int1132_t(x : std_logic_vector) return int1132_t;
subtype uint1133_t is unsigned(1132 downto 0);
constant uint1133_t_SLV_LEN : integer := 1133;
function uint1133_t_to_slv(x : uint1133_t) return std_logic_vector;
function slv_to_uint1133_t(x : std_logic_vector) return uint1133_t;
subtype int1133_t is signed(1132 downto 0);
constant int1133_t_SLV_LEN : integer := 1133;
function int1133_t_to_slv(x : int1133_t) return std_logic_vector;
function slv_to_int1133_t(x : std_logic_vector) return int1133_t;
subtype uint1134_t is unsigned(1133 downto 0);
constant uint1134_t_SLV_LEN : integer := 1134;
function uint1134_t_to_slv(x : uint1134_t) return std_logic_vector;
function slv_to_uint1134_t(x : std_logic_vector) return uint1134_t;
subtype int1134_t is signed(1133 downto 0);
constant int1134_t_SLV_LEN : integer := 1134;
function int1134_t_to_slv(x : int1134_t) return std_logic_vector;
function slv_to_int1134_t(x : std_logic_vector) return int1134_t;
subtype uint1135_t is unsigned(1134 downto 0);
constant uint1135_t_SLV_LEN : integer := 1135;
function uint1135_t_to_slv(x : uint1135_t) return std_logic_vector;
function slv_to_uint1135_t(x : std_logic_vector) return uint1135_t;
subtype int1135_t is signed(1134 downto 0);
constant int1135_t_SLV_LEN : integer := 1135;
function int1135_t_to_slv(x : int1135_t) return std_logic_vector;
function slv_to_int1135_t(x : std_logic_vector) return int1135_t;
subtype uint1136_t is unsigned(1135 downto 0);
constant uint1136_t_SLV_LEN : integer := 1136;
function uint1136_t_to_slv(x : uint1136_t) return std_logic_vector;
function slv_to_uint1136_t(x : std_logic_vector) return uint1136_t;
subtype int1136_t is signed(1135 downto 0);
constant int1136_t_SLV_LEN : integer := 1136;
function int1136_t_to_slv(x : int1136_t) return std_logic_vector;
function slv_to_int1136_t(x : std_logic_vector) return int1136_t;
subtype uint1137_t is unsigned(1136 downto 0);
constant uint1137_t_SLV_LEN : integer := 1137;
function uint1137_t_to_slv(x : uint1137_t) return std_logic_vector;
function slv_to_uint1137_t(x : std_logic_vector) return uint1137_t;
subtype int1137_t is signed(1136 downto 0);
constant int1137_t_SLV_LEN : integer := 1137;
function int1137_t_to_slv(x : int1137_t) return std_logic_vector;
function slv_to_int1137_t(x : std_logic_vector) return int1137_t;
subtype uint1138_t is unsigned(1137 downto 0);
constant uint1138_t_SLV_LEN : integer := 1138;
function uint1138_t_to_slv(x : uint1138_t) return std_logic_vector;
function slv_to_uint1138_t(x : std_logic_vector) return uint1138_t;
subtype int1138_t is signed(1137 downto 0);
constant int1138_t_SLV_LEN : integer := 1138;
function int1138_t_to_slv(x : int1138_t) return std_logic_vector;
function slv_to_int1138_t(x : std_logic_vector) return int1138_t;
subtype uint1139_t is unsigned(1138 downto 0);
constant uint1139_t_SLV_LEN : integer := 1139;
function uint1139_t_to_slv(x : uint1139_t) return std_logic_vector;
function slv_to_uint1139_t(x : std_logic_vector) return uint1139_t;
subtype int1139_t is signed(1138 downto 0);
constant int1139_t_SLV_LEN : integer := 1139;
function int1139_t_to_slv(x : int1139_t) return std_logic_vector;
function slv_to_int1139_t(x : std_logic_vector) return int1139_t;
subtype uint1140_t is unsigned(1139 downto 0);
constant uint1140_t_SLV_LEN : integer := 1140;
function uint1140_t_to_slv(x : uint1140_t) return std_logic_vector;
function slv_to_uint1140_t(x : std_logic_vector) return uint1140_t;
subtype int1140_t is signed(1139 downto 0);
constant int1140_t_SLV_LEN : integer := 1140;
function int1140_t_to_slv(x : int1140_t) return std_logic_vector;
function slv_to_int1140_t(x : std_logic_vector) return int1140_t;
subtype uint1141_t is unsigned(1140 downto 0);
constant uint1141_t_SLV_LEN : integer := 1141;
function uint1141_t_to_slv(x : uint1141_t) return std_logic_vector;
function slv_to_uint1141_t(x : std_logic_vector) return uint1141_t;
subtype int1141_t is signed(1140 downto 0);
constant int1141_t_SLV_LEN : integer := 1141;
function int1141_t_to_slv(x : int1141_t) return std_logic_vector;
function slv_to_int1141_t(x : std_logic_vector) return int1141_t;
subtype uint1142_t is unsigned(1141 downto 0);
constant uint1142_t_SLV_LEN : integer := 1142;
function uint1142_t_to_slv(x : uint1142_t) return std_logic_vector;
function slv_to_uint1142_t(x : std_logic_vector) return uint1142_t;
subtype int1142_t is signed(1141 downto 0);
constant int1142_t_SLV_LEN : integer := 1142;
function int1142_t_to_slv(x : int1142_t) return std_logic_vector;
function slv_to_int1142_t(x : std_logic_vector) return int1142_t;
subtype uint1143_t is unsigned(1142 downto 0);
constant uint1143_t_SLV_LEN : integer := 1143;
function uint1143_t_to_slv(x : uint1143_t) return std_logic_vector;
function slv_to_uint1143_t(x : std_logic_vector) return uint1143_t;
subtype int1143_t is signed(1142 downto 0);
constant int1143_t_SLV_LEN : integer := 1143;
function int1143_t_to_slv(x : int1143_t) return std_logic_vector;
function slv_to_int1143_t(x : std_logic_vector) return int1143_t;
subtype uint1144_t is unsigned(1143 downto 0);
constant uint1144_t_SLV_LEN : integer := 1144;
function uint1144_t_to_slv(x : uint1144_t) return std_logic_vector;
function slv_to_uint1144_t(x : std_logic_vector) return uint1144_t;
subtype int1144_t is signed(1143 downto 0);
constant int1144_t_SLV_LEN : integer := 1144;
function int1144_t_to_slv(x : int1144_t) return std_logic_vector;
function slv_to_int1144_t(x : std_logic_vector) return int1144_t;
subtype uint1145_t is unsigned(1144 downto 0);
constant uint1145_t_SLV_LEN : integer := 1145;
function uint1145_t_to_slv(x : uint1145_t) return std_logic_vector;
function slv_to_uint1145_t(x : std_logic_vector) return uint1145_t;
subtype int1145_t is signed(1144 downto 0);
constant int1145_t_SLV_LEN : integer := 1145;
function int1145_t_to_slv(x : int1145_t) return std_logic_vector;
function slv_to_int1145_t(x : std_logic_vector) return int1145_t;
subtype uint1146_t is unsigned(1145 downto 0);
constant uint1146_t_SLV_LEN : integer := 1146;
function uint1146_t_to_slv(x : uint1146_t) return std_logic_vector;
function slv_to_uint1146_t(x : std_logic_vector) return uint1146_t;
subtype int1146_t is signed(1145 downto 0);
constant int1146_t_SLV_LEN : integer := 1146;
function int1146_t_to_slv(x : int1146_t) return std_logic_vector;
function slv_to_int1146_t(x : std_logic_vector) return int1146_t;
subtype uint1147_t is unsigned(1146 downto 0);
constant uint1147_t_SLV_LEN : integer := 1147;
function uint1147_t_to_slv(x : uint1147_t) return std_logic_vector;
function slv_to_uint1147_t(x : std_logic_vector) return uint1147_t;
subtype int1147_t is signed(1146 downto 0);
constant int1147_t_SLV_LEN : integer := 1147;
function int1147_t_to_slv(x : int1147_t) return std_logic_vector;
function slv_to_int1147_t(x : std_logic_vector) return int1147_t;
subtype uint1148_t is unsigned(1147 downto 0);
constant uint1148_t_SLV_LEN : integer := 1148;
function uint1148_t_to_slv(x : uint1148_t) return std_logic_vector;
function slv_to_uint1148_t(x : std_logic_vector) return uint1148_t;
subtype int1148_t is signed(1147 downto 0);
constant int1148_t_SLV_LEN : integer := 1148;
function int1148_t_to_slv(x : int1148_t) return std_logic_vector;
function slv_to_int1148_t(x : std_logic_vector) return int1148_t;
subtype uint1149_t is unsigned(1148 downto 0);
constant uint1149_t_SLV_LEN : integer := 1149;
function uint1149_t_to_slv(x : uint1149_t) return std_logic_vector;
function slv_to_uint1149_t(x : std_logic_vector) return uint1149_t;
subtype int1149_t is signed(1148 downto 0);
constant int1149_t_SLV_LEN : integer := 1149;
function int1149_t_to_slv(x : int1149_t) return std_logic_vector;
function slv_to_int1149_t(x : std_logic_vector) return int1149_t;
subtype uint1150_t is unsigned(1149 downto 0);
constant uint1150_t_SLV_LEN : integer := 1150;
function uint1150_t_to_slv(x : uint1150_t) return std_logic_vector;
function slv_to_uint1150_t(x : std_logic_vector) return uint1150_t;
subtype int1150_t is signed(1149 downto 0);
constant int1150_t_SLV_LEN : integer := 1150;
function int1150_t_to_slv(x : int1150_t) return std_logic_vector;
function slv_to_int1150_t(x : std_logic_vector) return int1150_t;
subtype uint1151_t is unsigned(1150 downto 0);
constant uint1151_t_SLV_LEN : integer := 1151;
function uint1151_t_to_slv(x : uint1151_t) return std_logic_vector;
function slv_to_uint1151_t(x : std_logic_vector) return uint1151_t;
subtype int1151_t is signed(1150 downto 0);
constant int1151_t_SLV_LEN : integer := 1151;
function int1151_t_to_slv(x : int1151_t) return std_logic_vector;
function slv_to_int1151_t(x : std_logic_vector) return int1151_t;
subtype uint1152_t is unsigned(1151 downto 0);
constant uint1152_t_SLV_LEN : integer := 1152;
function uint1152_t_to_slv(x : uint1152_t) return std_logic_vector;
function slv_to_uint1152_t(x : std_logic_vector) return uint1152_t;
subtype int1152_t is signed(1151 downto 0);
constant int1152_t_SLV_LEN : integer := 1152;
function int1152_t_to_slv(x : int1152_t) return std_logic_vector;
function slv_to_int1152_t(x : std_logic_vector) return int1152_t;
subtype uint1153_t is unsigned(1152 downto 0);
constant uint1153_t_SLV_LEN : integer := 1153;
function uint1153_t_to_slv(x : uint1153_t) return std_logic_vector;
function slv_to_uint1153_t(x : std_logic_vector) return uint1153_t;
subtype int1153_t is signed(1152 downto 0);
constant int1153_t_SLV_LEN : integer := 1153;
function int1153_t_to_slv(x : int1153_t) return std_logic_vector;
function slv_to_int1153_t(x : std_logic_vector) return int1153_t;
subtype uint1154_t is unsigned(1153 downto 0);
constant uint1154_t_SLV_LEN : integer := 1154;
function uint1154_t_to_slv(x : uint1154_t) return std_logic_vector;
function slv_to_uint1154_t(x : std_logic_vector) return uint1154_t;
subtype int1154_t is signed(1153 downto 0);
constant int1154_t_SLV_LEN : integer := 1154;
function int1154_t_to_slv(x : int1154_t) return std_logic_vector;
function slv_to_int1154_t(x : std_logic_vector) return int1154_t;
subtype uint1155_t is unsigned(1154 downto 0);
constant uint1155_t_SLV_LEN : integer := 1155;
function uint1155_t_to_slv(x : uint1155_t) return std_logic_vector;
function slv_to_uint1155_t(x : std_logic_vector) return uint1155_t;
subtype int1155_t is signed(1154 downto 0);
constant int1155_t_SLV_LEN : integer := 1155;
function int1155_t_to_slv(x : int1155_t) return std_logic_vector;
function slv_to_int1155_t(x : std_logic_vector) return int1155_t;
subtype uint1156_t is unsigned(1155 downto 0);
constant uint1156_t_SLV_LEN : integer := 1156;
function uint1156_t_to_slv(x : uint1156_t) return std_logic_vector;
function slv_to_uint1156_t(x : std_logic_vector) return uint1156_t;
subtype int1156_t is signed(1155 downto 0);
constant int1156_t_SLV_LEN : integer := 1156;
function int1156_t_to_slv(x : int1156_t) return std_logic_vector;
function slv_to_int1156_t(x : std_logic_vector) return int1156_t;
subtype uint1157_t is unsigned(1156 downto 0);
constant uint1157_t_SLV_LEN : integer := 1157;
function uint1157_t_to_slv(x : uint1157_t) return std_logic_vector;
function slv_to_uint1157_t(x : std_logic_vector) return uint1157_t;
subtype int1157_t is signed(1156 downto 0);
constant int1157_t_SLV_LEN : integer := 1157;
function int1157_t_to_slv(x : int1157_t) return std_logic_vector;
function slv_to_int1157_t(x : std_logic_vector) return int1157_t;
subtype uint1158_t is unsigned(1157 downto 0);
constant uint1158_t_SLV_LEN : integer := 1158;
function uint1158_t_to_slv(x : uint1158_t) return std_logic_vector;
function slv_to_uint1158_t(x : std_logic_vector) return uint1158_t;
subtype int1158_t is signed(1157 downto 0);
constant int1158_t_SLV_LEN : integer := 1158;
function int1158_t_to_slv(x : int1158_t) return std_logic_vector;
function slv_to_int1158_t(x : std_logic_vector) return int1158_t;
subtype uint1159_t is unsigned(1158 downto 0);
constant uint1159_t_SLV_LEN : integer := 1159;
function uint1159_t_to_slv(x : uint1159_t) return std_logic_vector;
function slv_to_uint1159_t(x : std_logic_vector) return uint1159_t;
subtype int1159_t is signed(1158 downto 0);
constant int1159_t_SLV_LEN : integer := 1159;
function int1159_t_to_slv(x : int1159_t) return std_logic_vector;
function slv_to_int1159_t(x : std_logic_vector) return int1159_t;
subtype uint1160_t is unsigned(1159 downto 0);
constant uint1160_t_SLV_LEN : integer := 1160;
function uint1160_t_to_slv(x : uint1160_t) return std_logic_vector;
function slv_to_uint1160_t(x : std_logic_vector) return uint1160_t;
subtype int1160_t is signed(1159 downto 0);
constant int1160_t_SLV_LEN : integer := 1160;
function int1160_t_to_slv(x : int1160_t) return std_logic_vector;
function slv_to_int1160_t(x : std_logic_vector) return int1160_t;
subtype uint1161_t is unsigned(1160 downto 0);
constant uint1161_t_SLV_LEN : integer := 1161;
function uint1161_t_to_slv(x : uint1161_t) return std_logic_vector;
function slv_to_uint1161_t(x : std_logic_vector) return uint1161_t;
subtype int1161_t is signed(1160 downto 0);
constant int1161_t_SLV_LEN : integer := 1161;
function int1161_t_to_slv(x : int1161_t) return std_logic_vector;
function slv_to_int1161_t(x : std_logic_vector) return int1161_t;
subtype uint1162_t is unsigned(1161 downto 0);
constant uint1162_t_SLV_LEN : integer := 1162;
function uint1162_t_to_slv(x : uint1162_t) return std_logic_vector;
function slv_to_uint1162_t(x : std_logic_vector) return uint1162_t;
subtype int1162_t is signed(1161 downto 0);
constant int1162_t_SLV_LEN : integer := 1162;
function int1162_t_to_slv(x : int1162_t) return std_logic_vector;
function slv_to_int1162_t(x : std_logic_vector) return int1162_t;
subtype uint1163_t is unsigned(1162 downto 0);
constant uint1163_t_SLV_LEN : integer := 1163;
function uint1163_t_to_slv(x : uint1163_t) return std_logic_vector;
function slv_to_uint1163_t(x : std_logic_vector) return uint1163_t;
subtype int1163_t is signed(1162 downto 0);
constant int1163_t_SLV_LEN : integer := 1163;
function int1163_t_to_slv(x : int1163_t) return std_logic_vector;
function slv_to_int1163_t(x : std_logic_vector) return int1163_t;
subtype uint1164_t is unsigned(1163 downto 0);
constant uint1164_t_SLV_LEN : integer := 1164;
function uint1164_t_to_slv(x : uint1164_t) return std_logic_vector;
function slv_to_uint1164_t(x : std_logic_vector) return uint1164_t;
subtype int1164_t is signed(1163 downto 0);
constant int1164_t_SLV_LEN : integer := 1164;
function int1164_t_to_slv(x : int1164_t) return std_logic_vector;
function slv_to_int1164_t(x : std_logic_vector) return int1164_t;
subtype uint1165_t is unsigned(1164 downto 0);
constant uint1165_t_SLV_LEN : integer := 1165;
function uint1165_t_to_slv(x : uint1165_t) return std_logic_vector;
function slv_to_uint1165_t(x : std_logic_vector) return uint1165_t;
subtype int1165_t is signed(1164 downto 0);
constant int1165_t_SLV_LEN : integer := 1165;
function int1165_t_to_slv(x : int1165_t) return std_logic_vector;
function slv_to_int1165_t(x : std_logic_vector) return int1165_t;
subtype uint1166_t is unsigned(1165 downto 0);
constant uint1166_t_SLV_LEN : integer := 1166;
function uint1166_t_to_slv(x : uint1166_t) return std_logic_vector;
function slv_to_uint1166_t(x : std_logic_vector) return uint1166_t;
subtype int1166_t is signed(1165 downto 0);
constant int1166_t_SLV_LEN : integer := 1166;
function int1166_t_to_slv(x : int1166_t) return std_logic_vector;
function slv_to_int1166_t(x : std_logic_vector) return int1166_t;
subtype uint1167_t is unsigned(1166 downto 0);
constant uint1167_t_SLV_LEN : integer := 1167;
function uint1167_t_to_slv(x : uint1167_t) return std_logic_vector;
function slv_to_uint1167_t(x : std_logic_vector) return uint1167_t;
subtype int1167_t is signed(1166 downto 0);
constant int1167_t_SLV_LEN : integer := 1167;
function int1167_t_to_slv(x : int1167_t) return std_logic_vector;
function slv_to_int1167_t(x : std_logic_vector) return int1167_t;
subtype uint1168_t is unsigned(1167 downto 0);
constant uint1168_t_SLV_LEN : integer := 1168;
function uint1168_t_to_slv(x : uint1168_t) return std_logic_vector;
function slv_to_uint1168_t(x : std_logic_vector) return uint1168_t;
subtype int1168_t is signed(1167 downto 0);
constant int1168_t_SLV_LEN : integer := 1168;
function int1168_t_to_slv(x : int1168_t) return std_logic_vector;
function slv_to_int1168_t(x : std_logic_vector) return int1168_t;
subtype uint1169_t is unsigned(1168 downto 0);
constant uint1169_t_SLV_LEN : integer := 1169;
function uint1169_t_to_slv(x : uint1169_t) return std_logic_vector;
function slv_to_uint1169_t(x : std_logic_vector) return uint1169_t;
subtype int1169_t is signed(1168 downto 0);
constant int1169_t_SLV_LEN : integer := 1169;
function int1169_t_to_slv(x : int1169_t) return std_logic_vector;
function slv_to_int1169_t(x : std_logic_vector) return int1169_t;
subtype uint1170_t is unsigned(1169 downto 0);
constant uint1170_t_SLV_LEN : integer := 1170;
function uint1170_t_to_slv(x : uint1170_t) return std_logic_vector;
function slv_to_uint1170_t(x : std_logic_vector) return uint1170_t;
subtype int1170_t is signed(1169 downto 0);
constant int1170_t_SLV_LEN : integer := 1170;
function int1170_t_to_slv(x : int1170_t) return std_logic_vector;
function slv_to_int1170_t(x : std_logic_vector) return int1170_t;
subtype uint1171_t is unsigned(1170 downto 0);
constant uint1171_t_SLV_LEN : integer := 1171;
function uint1171_t_to_slv(x : uint1171_t) return std_logic_vector;
function slv_to_uint1171_t(x : std_logic_vector) return uint1171_t;
subtype int1171_t is signed(1170 downto 0);
constant int1171_t_SLV_LEN : integer := 1171;
function int1171_t_to_slv(x : int1171_t) return std_logic_vector;
function slv_to_int1171_t(x : std_logic_vector) return int1171_t;
subtype uint1172_t is unsigned(1171 downto 0);
constant uint1172_t_SLV_LEN : integer := 1172;
function uint1172_t_to_slv(x : uint1172_t) return std_logic_vector;
function slv_to_uint1172_t(x : std_logic_vector) return uint1172_t;
subtype int1172_t is signed(1171 downto 0);
constant int1172_t_SLV_LEN : integer := 1172;
function int1172_t_to_slv(x : int1172_t) return std_logic_vector;
function slv_to_int1172_t(x : std_logic_vector) return int1172_t;
subtype uint1173_t is unsigned(1172 downto 0);
constant uint1173_t_SLV_LEN : integer := 1173;
function uint1173_t_to_slv(x : uint1173_t) return std_logic_vector;
function slv_to_uint1173_t(x : std_logic_vector) return uint1173_t;
subtype int1173_t is signed(1172 downto 0);
constant int1173_t_SLV_LEN : integer := 1173;
function int1173_t_to_slv(x : int1173_t) return std_logic_vector;
function slv_to_int1173_t(x : std_logic_vector) return int1173_t;
subtype uint1174_t is unsigned(1173 downto 0);
constant uint1174_t_SLV_LEN : integer := 1174;
function uint1174_t_to_slv(x : uint1174_t) return std_logic_vector;
function slv_to_uint1174_t(x : std_logic_vector) return uint1174_t;
subtype int1174_t is signed(1173 downto 0);
constant int1174_t_SLV_LEN : integer := 1174;
function int1174_t_to_slv(x : int1174_t) return std_logic_vector;
function slv_to_int1174_t(x : std_logic_vector) return int1174_t;
subtype uint1175_t is unsigned(1174 downto 0);
constant uint1175_t_SLV_LEN : integer := 1175;
function uint1175_t_to_slv(x : uint1175_t) return std_logic_vector;
function slv_to_uint1175_t(x : std_logic_vector) return uint1175_t;
subtype int1175_t is signed(1174 downto 0);
constant int1175_t_SLV_LEN : integer := 1175;
function int1175_t_to_slv(x : int1175_t) return std_logic_vector;
function slv_to_int1175_t(x : std_logic_vector) return int1175_t;
subtype uint1176_t is unsigned(1175 downto 0);
constant uint1176_t_SLV_LEN : integer := 1176;
function uint1176_t_to_slv(x : uint1176_t) return std_logic_vector;
function slv_to_uint1176_t(x : std_logic_vector) return uint1176_t;
subtype int1176_t is signed(1175 downto 0);
constant int1176_t_SLV_LEN : integer := 1176;
function int1176_t_to_slv(x : int1176_t) return std_logic_vector;
function slv_to_int1176_t(x : std_logic_vector) return int1176_t;
subtype uint1177_t is unsigned(1176 downto 0);
constant uint1177_t_SLV_LEN : integer := 1177;
function uint1177_t_to_slv(x : uint1177_t) return std_logic_vector;
function slv_to_uint1177_t(x : std_logic_vector) return uint1177_t;
subtype int1177_t is signed(1176 downto 0);
constant int1177_t_SLV_LEN : integer := 1177;
function int1177_t_to_slv(x : int1177_t) return std_logic_vector;
function slv_to_int1177_t(x : std_logic_vector) return int1177_t;
subtype uint1178_t is unsigned(1177 downto 0);
constant uint1178_t_SLV_LEN : integer := 1178;
function uint1178_t_to_slv(x : uint1178_t) return std_logic_vector;
function slv_to_uint1178_t(x : std_logic_vector) return uint1178_t;
subtype int1178_t is signed(1177 downto 0);
constant int1178_t_SLV_LEN : integer := 1178;
function int1178_t_to_slv(x : int1178_t) return std_logic_vector;
function slv_to_int1178_t(x : std_logic_vector) return int1178_t;
subtype uint1179_t is unsigned(1178 downto 0);
constant uint1179_t_SLV_LEN : integer := 1179;
function uint1179_t_to_slv(x : uint1179_t) return std_logic_vector;
function slv_to_uint1179_t(x : std_logic_vector) return uint1179_t;
subtype int1179_t is signed(1178 downto 0);
constant int1179_t_SLV_LEN : integer := 1179;
function int1179_t_to_slv(x : int1179_t) return std_logic_vector;
function slv_to_int1179_t(x : std_logic_vector) return int1179_t;
subtype uint1180_t is unsigned(1179 downto 0);
constant uint1180_t_SLV_LEN : integer := 1180;
function uint1180_t_to_slv(x : uint1180_t) return std_logic_vector;
function slv_to_uint1180_t(x : std_logic_vector) return uint1180_t;
subtype int1180_t is signed(1179 downto 0);
constant int1180_t_SLV_LEN : integer := 1180;
function int1180_t_to_slv(x : int1180_t) return std_logic_vector;
function slv_to_int1180_t(x : std_logic_vector) return int1180_t;
subtype uint1181_t is unsigned(1180 downto 0);
constant uint1181_t_SLV_LEN : integer := 1181;
function uint1181_t_to_slv(x : uint1181_t) return std_logic_vector;
function slv_to_uint1181_t(x : std_logic_vector) return uint1181_t;
subtype int1181_t is signed(1180 downto 0);
constant int1181_t_SLV_LEN : integer := 1181;
function int1181_t_to_slv(x : int1181_t) return std_logic_vector;
function slv_to_int1181_t(x : std_logic_vector) return int1181_t;
subtype uint1182_t is unsigned(1181 downto 0);
constant uint1182_t_SLV_LEN : integer := 1182;
function uint1182_t_to_slv(x : uint1182_t) return std_logic_vector;
function slv_to_uint1182_t(x : std_logic_vector) return uint1182_t;
subtype int1182_t is signed(1181 downto 0);
constant int1182_t_SLV_LEN : integer := 1182;
function int1182_t_to_slv(x : int1182_t) return std_logic_vector;
function slv_to_int1182_t(x : std_logic_vector) return int1182_t;
subtype uint1183_t is unsigned(1182 downto 0);
constant uint1183_t_SLV_LEN : integer := 1183;
function uint1183_t_to_slv(x : uint1183_t) return std_logic_vector;
function slv_to_uint1183_t(x : std_logic_vector) return uint1183_t;
subtype int1183_t is signed(1182 downto 0);
constant int1183_t_SLV_LEN : integer := 1183;
function int1183_t_to_slv(x : int1183_t) return std_logic_vector;
function slv_to_int1183_t(x : std_logic_vector) return int1183_t;
subtype uint1184_t is unsigned(1183 downto 0);
constant uint1184_t_SLV_LEN : integer := 1184;
function uint1184_t_to_slv(x : uint1184_t) return std_logic_vector;
function slv_to_uint1184_t(x : std_logic_vector) return uint1184_t;
subtype int1184_t is signed(1183 downto 0);
constant int1184_t_SLV_LEN : integer := 1184;
function int1184_t_to_slv(x : int1184_t) return std_logic_vector;
function slv_to_int1184_t(x : std_logic_vector) return int1184_t;
subtype uint1185_t is unsigned(1184 downto 0);
constant uint1185_t_SLV_LEN : integer := 1185;
function uint1185_t_to_slv(x : uint1185_t) return std_logic_vector;
function slv_to_uint1185_t(x : std_logic_vector) return uint1185_t;
subtype int1185_t is signed(1184 downto 0);
constant int1185_t_SLV_LEN : integer := 1185;
function int1185_t_to_slv(x : int1185_t) return std_logic_vector;
function slv_to_int1185_t(x : std_logic_vector) return int1185_t;
subtype uint1186_t is unsigned(1185 downto 0);
constant uint1186_t_SLV_LEN : integer := 1186;
function uint1186_t_to_slv(x : uint1186_t) return std_logic_vector;
function slv_to_uint1186_t(x : std_logic_vector) return uint1186_t;
subtype int1186_t is signed(1185 downto 0);
constant int1186_t_SLV_LEN : integer := 1186;
function int1186_t_to_slv(x : int1186_t) return std_logic_vector;
function slv_to_int1186_t(x : std_logic_vector) return int1186_t;
subtype uint1187_t is unsigned(1186 downto 0);
constant uint1187_t_SLV_LEN : integer := 1187;
function uint1187_t_to_slv(x : uint1187_t) return std_logic_vector;
function slv_to_uint1187_t(x : std_logic_vector) return uint1187_t;
subtype int1187_t is signed(1186 downto 0);
constant int1187_t_SLV_LEN : integer := 1187;
function int1187_t_to_slv(x : int1187_t) return std_logic_vector;
function slv_to_int1187_t(x : std_logic_vector) return int1187_t;
subtype uint1188_t is unsigned(1187 downto 0);
constant uint1188_t_SLV_LEN : integer := 1188;
function uint1188_t_to_slv(x : uint1188_t) return std_logic_vector;
function slv_to_uint1188_t(x : std_logic_vector) return uint1188_t;
subtype int1188_t is signed(1187 downto 0);
constant int1188_t_SLV_LEN : integer := 1188;
function int1188_t_to_slv(x : int1188_t) return std_logic_vector;
function slv_to_int1188_t(x : std_logic_vector) return int1188_t;
subtype uint1189_t is unsigned(1188 downto 0);
constant uint1189_t_SLV_LEN : integer := 1189;
function uint1189_t_to_slv(x : uint1189_t) return std_logic_vector;
function slv_to_uint1189_t(x : std_logic_vector) return uint1189_t;
subtype int1189_t is signed(1188 downto 0);
constant int1189_t_SLV_LEN : integer := 1189;
function int1189_t_to_slv(x : int1189_t) return std_logic_vector;
function slv_to_int1189_t(x : std_logic_vector) return int1189_t;
subtype uint1190_t is unsigned(1189 downto 0);
constant uint1190_t_SLV_LEN : integer := 1190;
function uint1190_t_to_slv(x : uint1190_t) return std_logic_vector;
function slv_to_uint1190_t(x : std_logic_vector) return uint1190_t;
subtype int1190_t is signed(1189 downto 0);
constant int1190_t_SLV_LEN : integer := 1190;
function int1190_t_to_slv(x : int1190_t) return std_logic_vector;
function slv_to_int1190_t(x : std_logic_vector) return int1190_t;
subtype uint1191_t is unsigned(1190 downto 0);
constant uint1191_t_SLV_LEN : integer := 1191;
function uint1191_t_to_slv(x : uint1191_t) return std_logic_vector;
function slv_to_uint1191_t(x : std_logic_vector) return uint1191_t;
subtype int1191_t is signed(1190 downto 0);
constant int1191_t_SLV_LEN : integer := 1191;
function int1191_t_to_slv(x : int1191_t) return std_logic_vector;
function slv_to_int1191_t(x : std_logic_vector) return int1191_t;
subtype uint1192_t is unsigned(1191 downto 0);
constant uint1192_t_SLV_LEN : integer := 1192;
function uint1192_t_to_slv(x : uint1192_t) return std_logic_vector;
function slv_to_uint1192_t(x : std_logic_vector) return uint1192_t;
subtype int1192_t is signed(1191 downto 0);
constant int1192_t_SLV_LEN : integer := 1192;
function int1192_t_to_slv(x : int1192_t) return std_logic_vector;
function slv_to_int1192_t(x : std_logic_vector) return int1192_t;
subtype uint1193_t is unsigned(1192 downto 0);
constant uint1193_t_SLV_LEN : integer := 1193;
function uint1193_t_to_slv(x : uint1193_t) return std_logic_vector;
function slv_to_uint1193_t(x : std_logic_vector) return uint1193_t;
subtype int1193_t is signed(1192 downto 0);
constant int1193_t_SLV_LEN : integer := 1193;
function int1193_t_to_slv(x : int1193_t) return std_logic_vector;
function slv_to_int1193_t(x : std_logic_vector) return int1193_t;
subtype uint1194_t is unsigned(1193 downto 0);
constant uint1194_t_SLV_LEN : integer := 1194;
function uint1194_t_to_slv(x : uint1194_t) return std_logic_vector;
function slv_to_uint1194_t(x : std_logic_vector) return uint1194_t;
subtype int1194_t is signed(1193 downto 0);
constant int1194_t_SLV_LEN : integer := 1194;
function int1194_t_to_slv(x : int1194_t) return std_logic_vector;
function slv_to_int1194_t(x : std_logic_vector) return int1194_t;
subtype uint1195_t is unsigned(1194 downto 0);
constant uint1195_t_SLV_LEN : integer := 1195;
function uint1195_t_to_slv(x : uint1195_t) return std_logic_vector;
function slv_to_uint1195_t(x : std_logic_vector) return uint1195_t;
subtype int1195_t is signed(1194 downto 0);
constant int1195_t_SLV_LEN : integer := 1195;
function int1195_t_to_slv(x : int1195_t) return std_logic_vector;
function slv_to_int1195_t(x : std_logic_vector) return int1195_t;
subtype uint1196_t is unsigned(1195 downto 0);
constant uint1196_t_SLV_LEN : integer := 1196;
function uint1196_t_to_slv(x : uint1196_t) return std_logic_vector;
function slv_to_uint1196_t(x : std_logic_vector) return uint1196_t;
subtype int1196_t is signed(1195 downto 0);
constant int1196_t_SLV_LEN : integer := 1196;
function int1196_t_to_slv(x : int1196_t) return std_logic_vector;
function slv_to_int1196_t(x : std_logic_vector) return int1196_t;
subtype uint1197_t is unsigned(1196 downto 0);
constant uint1197_t_SLV_LEN : integer := 1197;
function uint1197_t_to_slv(x : uint1197_t) return std_logic_vector;
function slv_to_uint1197_t(x : std_logic_vector) return uint1197_t;
subtype int1197_t is signed(1196 downto 0);
constant int1197_t_SLV_LEN : integer := 1197;
function int1197_t_to_slv(x : int1197_t) return std_logic_vector;
function slv_to_int1197_t(x : std_logic_vector) return int1197_t;
subtype uint1198_t is unsigned(1197 downto 0);
constant uint1198_t_SLV_LEN : integer := 1198;
function uint1198_t_to_slv(x : uint1198_t) return std_logic_vector;
function slv_to_uint1198_t(x : std_logic_vector) return uint1198_t;
subtype int1198_t is signed(1197 downto 0);
constant int1198_t_SLV_LEN : integer := 1198;
function int1198_t_to_slv(x : int1198_t) return std_logic_vector;
function slv_to_int1198_t(x : std_logic_vector) return int1198_t;
subtype uint1199_t is unsigned(1198 downto 0);
constant uint1199_t_SLV_LEN : integer := 1199;
function uint1199_t_to_slv(x : uint1199_t) return std_logic_vector;
function slv_to_uint1199_t(x : std_logic_vector) return uint1199_t;
subtype int1199_t is signed(1198 downto 0);
constant int1199_t_SLV_LEN : integer := 1199;
function int1199_t_to_slv(x : int1199_t) return std_logic_vector;
function slv_to_int1199_t(x : std_logic_vector) return int1199_t;
subtype uint1200_t is unsigned(1199 downto 0);
constant uint1200_t_SLV_LEN : integer := 1200;
function uint1200_t_to_slv(x : uint1200_t) return std_logic_vector;
function slv_to_uint1200_t(x : std_logic_vector) return uint1200_t;
subtype int1200_t is signed(1199 downto 0);
constant int1200_t_SLV_LEN : integer := 1200;
function int1200_t_to_slv(x : int1200_t) return std_logic_vector;
function slv_to_int1200_t(x : std_logic_vector) return int1200_t;
subtype uint1201_t is unsigned(1200 downto 0);
constant uint1201_t_SLV_LEN : integer := 1201;
function uint1201_t_to_slv(x : uint1201_t) return std_logic_vector;
function slv_to_uint1201_t(x : std_logic_vector) return uint1201_t;
subtype int1201_t is signed(1200 downto 0);
constant int1201_t_SLV_LEN : integer := 1201;
function int1201_t_to_slv(x : int1201_t) return std_logic_vector;
function slv_to_int1201_t(x : std_logic_vector) return int1201_t;
subtype uint1202_t is unsigned(1201 downto 0);
constant uint1202_t_SLV_LEN : integer := 1202;
function uint1202_t_to_slv(x : uint1202_t) return std_logic_vector;
function slv_to_uint1202_t(x : std_logic_vector) return uint1202_t;
subtype int1202_t is signed(1201 downto 0);
constant int1202_t_SLV_LEN : integer := 1202;
function int1202_t_to_slv(x : int1202_t) return std_logic_vector;
function slv_to_int1202_t(x : std_logic_vector) return int1202_t;
subtype uint1203_t is unsigned(1202 downto 0);
constant uint1203_t_SLV_LEN : integer := 1203;
function uint1203_t_to_slv(x : uint1203_t) return std_logic_vector;
function slv_to_uint1203_t(x : std_logic_vector) return uint1203_t;
subtype int1203_t is signed(1202 downto 0);
constant int1203_t_SLV_LEN : integer := 1203;
function int1203_t_to_slv(x : int1203_t) return std_logic_vector;
function slv_to_int1203_t(x : std_logic_vector) return int1203_t;
subtype uint1204_t is unsigned(1203 downto 0);
constant uint1204_t_SLV_LEN : integer := 1204;
function uint1204_t_to_slv(x : uint1204_t) return std_logic_vector;
function slv_to_uint1204_t(x : std_logic_vector) return uint1204_t;
subtype int1204_t is signed(1203 downto 0);
constant int1204_t_SLV_LEN : integer := 1204;
function int1204_t_to_slv(x : int1204_t) return std_logic_vector;
function slv_to_int1204_t(x : std_logic_vector) return int1204_t;
subtype uint1205_t is unsigned(1204 downto 0);
constant uint1205_t_SLV_LEN : integer := 1205;
function uint1205_t_to_slv(x : uint1205_t) return std_logic_vector;
function slv_to_uint1205_t(x : std_logic_vector) return uint1205_t;
subtype int1205_t is signed(1204 downto 0);
constant int1205_t_SLV_LEN : integer := 1205;
function int1205_t_to_slv(x : int1205_t) return std_logic_vector;
function slv_to_int1205_t(x : std_logic_vector) return int1205_t;
subtype uint1206_t is unsigned(1205 downto 0);
constant uint1206_t_SLV_LEN : integer := 1206;
function uint1206_t_to_slv(x : uint1206_t) return std_logic_vector;
function slv_to_uint1206_t(x : std_logic_vector) return uint1206_t;
subtype int1206_t is signed(1205 downto 0);
constant int1206_t_SLV_LEN : integer := 1206;
function int1206_t_to_slv(x : int1206_t) return std_logic_vector;
function slv_to_int1206_t(x : std_logic_vector) return int1206_t;
subtype uint1207_t is unsigned(1206 downto 0);
constant uint1207_t_SLV_LEN : integer := 1207;
function uint1207_t_to_slv(x : uint1207_t) return std_logic_vector;
function slv_to_uint1207_t(x : std_logic_vector) return uint1207_t;
subtype int1207_t is signed(1206 downto 0);
constant int1207_t_SLV_LEN : integer := 1207;
function int1207_t_to_slv(x : int1207_t) return std_logic_vector;
function slv_to_int1207_t(x : std_logic_vector) return int1207_t;
subtype uint1208_t is unsigned(1207 downto 0);
constant uint1208_t_SLV_LEN : integer := 1208;
function uint1208_t_to_slv(x : uint1208_t) return std_logic_vector;
function slv_to_uint1208_t(x : std_logic_vector) return uint1208_t;
subtype int1208_t is signed(1207 downto 0);
constant int1208_t_SLV_LEN : integer := 1208;
function int1208_t_to_slv(x : int1208_t) return std_logic_vector;
function slv_to_int1208_t(x : std_logic_vector) return int1208_t;
subtype uint1209_t is unsigned(1208 downto 0);
constant uint1209_t_SLV_LEN : integer := 1209;
function uint1209_t_to_slv(x : uint1209_t) return std_logic_vector;
function slv_to_uint1209_t(x : std_logic_vector) return uint1209_t;
subtype int1209_t is signed(1208 downto 0);
constant int1209_t_SLV_LEN : integer := 1209;
function int1209_t_to_slv(x : int1209_t) return std_logic_vector;
function slv_to_int1209_t(x : std_logic_vector) return int1209_t;
subtype uint1210_t is unsigned(1209 downto 0);
constant uint1210_t_SLV_LEN : integer := 1210;
function uint1210_t_to_slv(x : uint1210_t) return std_logic_vector;
function slv_to_uint1210_t(x : std_logic_vector) return uint1210_t;
subtype int1210_t is signed(1209 downto 0);
constant int1210_t_SLV_LEN : integer := 1210;
function int1210_t_to_slv(x : int1210_t) return std_logic_vector;
function slv_to_int1210_t(x : std_logic_vector) return int1210_t;
subtype uint1211_t is unsigned(1210 downto 0);
constant uint1211_t_SLV_LEN : integer := 1211;
function uint1211_t_to_slv(x : uint1211_t) return std_logic_vector;
function slv_to_uint1211_t(x : std_logic_vector) return uint1211_t;
subtype int1211_t is signed(1210 downto 0);
constant int1211_t_SLV_LEN : integer := 1211;
function int1211_t_to_slv(x : int1211_t) return std_logic_vector;
function slv_to_int1211_t(x : std_logic_vector) return int1211_t;
subtype uint1212_t is unsigned(1211 downto 0);
constant uint1212_t_SLV_LEN : integer := 1212;
function uint1212_t_to_slv(x : uint1212_t) return std_logic_vector;
function slv_to_uint1212_t(x : std_logic_vector) return uint1212_t;
subtype int1212_t is signed(1211 downto 0);
constant int1212_t_SLV_LEN : integer := 1212;
function int1212_t_to_slv(x : int1212_t) return std_logic_vector;
function slv_to_int1212_t(x : std_logic_vector) return int1212_t;
subtype uint1213_t is unsigned(1212 downto 0);
constant uint1213_t_SLV_LEN : integer := 1213;
function uint1213_t_to_slv(x : uint1213_t) return std_logic_vector;
function slv_to_uint1213_t(x : std_logic_vector) return uint1213_t;
subtype int1213_t is signed(1212 downto 0);
constant int1213_t_SLV_LEN : integer := 1213;
function int1213_t_to_slv(x : int1213_t) return std_logic_vector;
function slv_to_int1213_t(x : std_logic_vector) return int1213_t;
subtype uint1214_t is unsigned(1213 downto 0);
constant uint1214_t_SLV_LEN : integer := 1214;
function uint1214_t_to_slv(x : uint1214_t) return std_logic_vector;
function slv_to_uint1214_t(x : std_logic_vector) return uint1214_t;
subtype int1214_t is signed(1213 downto 0);
constant int1214_t_SLV_LEN : integer := 1214;
function int1214_t_to_slv(x : int1214_t) return std_logic_vector;
function slv_to_int1214_t(x : std_logic_vector) return int1214_t;
subtype uint1215_t is unsigned(1214 downto 0);
constant uint1215_t_SLV_LEN : integer := 1215;
function uint1215_t_to_slv(x : uint1215_t) return std_logic_vector;
function slv_to_uint1215_t(x : std_logic_vector) return uint1215_t;
subtype int1215_t is signed(1214 downto 0);
constant int1215_t_SLV_LEN : integer := 1215;
function int1215_t_to_slv(x : int1215_t) return std_logic_vector;
function slv_to_int1215_t(x : std_logic_vector) return int1215_t;
subtype uint1216_t is unsigned(1215 downto 0);
constant uint1216_t_SLV_LEN : integer := 1216;
function uint1216_t_to_slv(x : uint1216_t) return std_logic_vector;
function slv_to_uint1216_t(x : std_logic_vector) return uint1216_t;
subtype int1216_t is signed(1215 downto 0);
constant int1216_t_SLV_LEN : integer := 1216;
function int1216_t_to_slv(x : int1216_t) return std_logic_vector;
function slv_to_int1216_t(x : std_logic_vector) return int1216_t;
subtype uint1217_t is unsigned(1216 downto 0);
constant uint1217_t_SLV_LEN : integer := 1217;
function uint1217_t_to_slv(x : uint1217_t) return std_logic_vector;
function slv_to_uint1217_t(x : std_logic_vector) return uint1217_t;
subtype int1217_t is signed(1216 downto 0);
constant int1217_t_SLV_LEN : integer := 1217;
function int1217_t_to_slv(x : int1217_t) return std_logic_vector;
function slv_to_int1217_t(x : std_logic_vector) return int1217_t;
subtype uint1218_t is unsigned(1217 downto 0);
constant uint1218_t_SLV_LEN : integer := 1218;
function uint1218_t_to_slv(x : uint1218_t) return std_logic_vector;
function slv_to_uint1218_t(x : std_logic_vector) return uint1218_t;
subtype int1218_t is signed(1217 downto 0);
constant int1218_t_SLV_LEN : integer := 1218;
function int1218_t_to_slv(x : int1218_t) return std_logic_vector;
function slv_to_int1218_t(x : std_logic_vector) return int1218_t;
subtype uint1219_t is unsigned(1218 downto 0);
constant uint1219_t_SLV_LEN : integer := 1219;
function uint1219_t_to_slv(x : uint1219_t) return std_logic_vector;
function slv_to_uint1219_t(x : std_logic_vector) return uint1219_t;
subtype int1219_t is signed(1218 downto 0);
constant int1219_t_SLV_LEN : integer := 1219;
function int1219_t_to_slv(x : int1219_t) return std_logic_vector;
function slv_to_int1219_t(x : std_logic_vector) return int1219_t;
subtype uint1220_t is unsigned(1219 downto 0);
constant uint1220_t_SLV_LEN : integer := 1220;
function uint1220_t_to_slv(x : uint1220_t) return std_logic_vector;
function slv_to_uint1220_t(x : std_logic_vector) return uint1220_t;
subtype int1220_t is signed(1219 downto 0);
constant int1220_t_SLV_LEN : integer := 1220;
function int1220_t_to_slv(x : int1220_t) return std_logic_vector;
function slv_to_int1220_t(x : std_logic_vector) return int1220_t;
subtype uint1221_t is unsigned(1220 downto 0);
constant uint1221_t_SLV_LEN : integer := 1221;
function uint1221_t_to_slv(x : uint1221_t) return std_logic_vector;
function slv_to_uint1221_t(x : std_logic_vector) return uint1221_t;
subtype int1221_t is signed(1220 downto 0);
constant int1221_t_SLV_LEN : integer := 1221;
function int1221_t_to_slv(x : int1221_t) return std_logic_vector;
function slv_to_int1221_t(x : std_logic_vector) return int1221_t;
subtype uint1222_t is unsigned(1221 downto 0);
constant uint1222_t_SLV_LEN : integer := 1222;
function uint1222_t_to_slv(x : uint1222_t) return std_logic_vector;
function slv_to_uint1222_t(x : std_logic_vector) return uint1222_t;
subtype int1222_t is signed(1221 downto 0);
constant int1222_t_SLV_LEN : integer := 1222;
function int1222_t_to_slv(x : int1222_t) return std_logic_vector;
function slv_to_int1222_t(x : std_logic_vector) return int1222_t;
subtype uint1223_t is unsigned(1222 downto 0);
constant uint1223_t_SLV_LEN : integer := 1223;
function uint1223_t_to_slv(x : uint1223_t) return std_logic_vector;
function slv_to_uint1223_t(x : std_logic_vector) return uint1223_t;
subtype int1223_t is signed(1222 downto 0);
constant int1223_t_SLV_LEN : integer := 1223;
function int1223_t_to_slv(x : int1223_t) return std_logic_vector;
function slv_to_int1223_t(x : std_logic_vector) return int1223_t;
subtype uint1224_t is unsigned(1223 downto 0);
constant uint1224_t_SLV_LEN : integer := 1224;
function uint1224_t_to_slv(x : uint1224_t) return std_logic_vector;
function slv_to_uint1224_t(x : std_logic_vector) return uint1224_t;
subtype int1224_t is signed(1223 downto 0);
constant int1224_t_SLV_LEN : integer := 1224;
function int1224_t_to_slv(x : int1224_t) return std_logic_vector;
function slv_to_int1224_t(x : std_logic_vector) return int1224_t;
subtype uint1225_t is unsigned(1224 downto 0);
constant uint1225_t_SLV_LEN : integer := 1225;
function uint1225_t_to_slv(x : uint1225_t) return std_logic_vector;
function slv_to_uint1225_t(x : std_logic_vector) return uint1225_t;
subtype int1225_t is signed(1224 downto 0);
constant int1225_t_SLV_LEN : integer := 1225;
function int1225_t_to_slv(x : int1225_t) return std_logic_vector;
function slv_to_int1225_t(x : std_logic_vector) return int1225_t;
subtype uint1226_t is unsigned(1225 downto 0);
constant uint1226_t_SLV_LEN : integer := 1226;
function uint1226_t_to_slv(x : uint1226_t) return std_logic_vector;
function slv_to_uint1226_t(x : std_logic_vector) return uint1226_t;
subtype int1226_t is signed(1225 downto 0);
constant int1226_t_SLV_LEN : integer := 1226;
function int1226_t_to_slv(x : int1226_t) return std_logic_vector;
function slv_to_int1226_t(x : std_logic_vector) return int1226_t;
subtype uint1227_t is unsigned(1226 downto 0);
constant uint1227_t_SLV_LEN : integer := 1227;
function uint1227_t_to_slv(x : uint1227_t) return std_logic_vector;
function slv_to_uint1227_t(x : std_logic_vector) return uint1227_t;
subtype int1227_t is signed(1226 downto 0);
constant int1227_t_SLV_LEN : integer := 1227;
function int1227_t_to_slv(x : int1227_t) return std_logic_vector;
function slv_to_int1227_t(x : std_logic_vector) return int1227_t;
subtype uint1228_t is unsigned(1227 downto 0);
constant uint1228_t_SLV_LEN : integer := 1228;
function uint1228_t_to_slv(x : uint1228_t) return std_logic_vector;
function slv_to_uint1228_t(x : std_logic_vector) return uint1228_t;
subtype int1228_t is signed(1227 downto 0);
constant int1228_t_SLV_LEN : integer := 1228;
function int1228_t_to_slv(x : int1228_t) return std_logic_vector;
function slv_to_int1228_t(x : std_logic_vector) return int1228_t;
subtype uint1229_t is unsigned(1228 downto 0);
constant uint1229_t_SLV_LEN : integer := 1229;
function uint1229_t_to_slv(x : uint1229_t) return std_logic_vector;
function slv_to_uint1229_t(x : std_logic_vector) return uint1229_t;
subtype int1229_t is signed(1228 downto 0);
constant int1229_t_SLV_LEN : integer := 1229;
function int1229_t_to_slv(x : int1229_t) return std_logic_vector;
function slv_to_int1229_t(x : std_logic_vector) return int1229_t;
subtype uint1230_t is unsigned(1229 downto 0);
constant uint1230_t_SLV_LEN : integer := 1230;
function uint1230_t_to_slv(x : uint1230_t) return std_logic_vector;
function slv_to_uint1230_t(x : std_logic_vector) return uint1230_t;
subtype int1230_t is signed(1229 downto 0);
constant int1230_t_SLV_LEN : integer := 1230;
function int1230_t_to_slv(x : int1230_t) return std_logic_vector;
function slv_to_int1230_t(x : std_logic_vector) return int1230_t;
subtype uint1231_t is unsigned(1230 downto 0);
constant uint1231_t_SLV_LEN : integer := 1231;
function uint1231_t_to_slv(x : uint1231_t) return std_logic_vector;
function slv_to_uint1231_t(x : std_logic_vector) return uint1231_t;
subtype int1231_t is signed(1230 downto 0);
constant int1231_t_SLV_LEN : integer := 1231;
function int1231_t_to_slv(x : int1231_t) return std_logic_vector;
function slv_to_int1231_t(x : std_logic_vector) return int1231_t;
subtype uint1232_t is unsigned(1231 downto 0);
constant uint1232_t_SLV_LEN : integer := 1232;
function uint1232_t_to_slv(x : uint1232_t) return std_logic_vector;
function slv_to_uint1232_t(x : std_logic_vector) return uint1232_t;
subtype int1232_t is signed(1231 downto 0);
constant int1232_t_SLV_LEN : integer := 1232;
function int1232_t_to_slv(x : int1232_t) return std_logic_vector;
function slv_to_int1232_t(x : std_logic_vector) return int1232_t;
subtype uint1233_t is unsigned(1232 downto 0);
constant uint1233_t_SLV_LEN : integer := 1233;
function uint1233_t_to_slv(x : uint1233_t) return std_logic_vector;
function slv_to_uint1233_t(x : std_logic_vector) return uint1233_t;
subtype int1233_t is signed(1232 downto 0);
constant int1233_t_SLV_LEN : integer := 1233;
function int1233_t_to_slv(x : int1233_t) return std_logic_vector;
function slv_to_int1233_t(x : std_logic_vector) return int1233_t;
subtype uint1234_t is unsigned(1233 downto 0);
constant uint1234_t_SLV_LEN : integer := 1234;
function uint1234_t_to_slv(x : uint1234_t) return std_logic_vector;
function slv_to_uint1234_t(x : std_logic_vector) return uint1234_t;
subtype int1234_t is signed(1233 downto 0);
constant int1234_t_SLV_LEN : integer := 1234;
function int1234_t_to_slv(x : int1234_t) return std_logic_vector;
function slv_to_int1234_t(x : std_logic_vector) return int1234_t;
subtype uint1235_t is unsigned(1234 downto 0);
constant uint1235_t_SLV_LEN : integer := 1235;
function uint1235_t_to_slv(x : uint1235_t) return std_logic_vector;
function slv_to_uint1235_t(x : std_logic_vector) return uint1235_t;
subtype int1235_t is signed(1234 downto 0);
constant int1235_t_SLV_LEN : integer := 1235;
function int1235_t_to_slv(x : int1235_t) return std_logic_vector;
function slv_to_int1235_t(x : std_logic_vector) return int1235_t;
subtype uint1236_t is unsigned(1235 downto 0);
constant uint1236_t_SLV_LEN : integer := 1236;
function uint1236_t_to_slv(x : uint1236_t) return std_logic_vector;
function slv_to_uint1236_t(x : std_logic_vector) return uint1236_t;
subtype int1236_t is signed(1235 downto 0);
constant int1236_t_SLV_LEN : integer := 1236;
function int1236_t_to_slv(x : int1236_t) return std_logic_vector;
function slv_to_int1236_t(x : std_logic_vector) return int1236_t;
subtype uint1237_t is unsigned(1236 downto 0);
constant uint1237_t_SLV_LEN : integer := 1237;
function uint1237_t_to_slv(x : uint1237_t) return std_logic_vector;
function slv_to_uint1237_t(x : std_logic_vector) return uint1237_t;
subtype int1237_t is signed(1236 downto 0);
constant int1237_t_SLV_LEN : integer := 1237;
function int1237_t_to_slv(x : int1237_t) return std_logic_vector;
function slv_to_int1237_t(x : std_logic_vector) return int1237_t;
subtype uint1238_t is unsigned(1237 downto 0);
constant uint1238_t_SLV_LEN : integer := 1238;
function uint1238_t_to_slv(x : uint1238_t) return std_logic_vector;
function slv_to_uint1238_t(x : std_logic_vector) return uint1238_t;
subtype int1238_t is signed(1237 downto 0);
constant int1238_t_SLV_LEN : integer := 1238;
function int1238_t_to_slv(x : int1238_t) return std_logic_vector;
function slv_to_int1238_t(x : std_logic_vector) return int1238_t;
subtype uint1239_t is unsigned(1238 downto 0);
constant uint1239_t_SLV_LEN : integer := 1239;
function uint1239_t_to_slv(x : uint1239_t) return std_logic_vector;
function slv_to_uint1239_t(x : std_logic_vector) return uint1239_t;
subtype int1239_t is signed(1238 downto 0);
constant int1239_t_SLV_LEN : integer := 1239;
function int1239_t_to_slv(x : int1239_t) return std_logic_vector;
function slv_to_int1239_t(x : std_logic_vector) return int1239_t;
subtype uint1240_t is unsigned(1239 downto 0);
constant uint1240_t_SLV_LEN : integer := 1240;
function uint1240_t_to_slv(x : uint1240_t) return std_logic_vector;
function slv_to_uint1240_t(x : std_logic_vector) return uint1240_t;
subtype int1240_t is signed(1239 downto 0);
constant int1240_t_SLV_LEN : integer := 1240;
function int1240_t_to_slv(x : int1240_t) return std_logic_vector;
function slv_to_int1240_t(x : std_logic_vector) return int1240_t;
subtype uint1241_t is unsigned(1240 downto 0);
constant uint1241_t_SLV_LEN : integer := 1241;
function uint1241_t_to_slv(x : uint1241_t) return std_logic_vector;
function slv_to_uint1241_t(x : std_logic_vector) return uint1241_t;
subtype int1241_t is signed(1240 downto 0);
constant int1241_t_SLV_LEN : integer := 1241;
function int1241_t_to_slv(x : int1241_t) return std_logic_vector;
function slv_to_int1241_t(x : std_logic_vector) return int1241_t;
subtype uint1242_t is unsigned(1241 downto 0);
constant uint1242_t_SLV_LEN : integer := 1242;
function uint1242_t_to_slv(x : uint1242_t) return std_logic_vector;
function slv_to_uint1242_t(x : std_logic_vector) return uint1242_t;
subtype int1242_t is signed(1241 downto 0);
constant int1242_t_SLV_LEN : integer := 1242;
function int1242_t_to_slv(x : int1242_t) return std_logic_vector;
function slv_to_int1242_t(x : std_logic_vector) return int1242_t;
subtype uint1243_t is unsigned(1242 downto 0);
constant uint1243_t_SLV_LEN : integer := 1243;
function uint1243_t_to_slv(x : uint1243_t) return std_logic_vector;
function slv_to_uint1243_t(x : std_logic_vector) return uint1243_t;
subtype int1243_t is signed(1242 downto 0);
constant int1243_t_SLV_LEN : integer := 1243;
function int1243_t_to_slv(x : int1243_t) return std_logic_vector;
function slv_to_int1243_t(x : std_logic_vector) return int1243_t;
subtype uint1244_t is unsigned(1243 downto 0);
constant uint1244_t_SLV_LEN : integer := 1244;
function uint1244_t_to_slv(x : uint1244_t) return std_logic_vector;
function slv_to_uint1244_t(x : std_logic_vector) return uint1244_t;
subtype int1244_t is signed(1243 downto 0);
constant int1244_t_SLV_LEN : integer := 1244;
function int1244_t_to_slv(x : int1244_t) return std_logic_vector;
function slv_to_int1244_t(x : std_logic_vector) return int1244_t;
subtype uint1245_t is unsigned(1244 downto 0);
constant uint1245_t_SLV_LEN : integer := 1245;
function uint1245_t_to_slv(x : uint1245_t) return std_logic_vector;
function slv_to_uint1245_t(x : std_logic_vector) return uint1245_t;
subtype int1245_t is signed(1244 downto 0);
constant int1245_t_SLV_LEN : integer := 1245;
function int1245_t_to_slv(x : int1245_t) return std_logic_vector;
function slv_to_int1245_t(x : std_logic_vector) return int1245_t;
subtype uint1246_t is unsigned(1245 downto 0);
constant uint1246_t_SLV_LEN : integer := 1246;
function uint1246_t_to_slv(x : uint1246_t) return std_logic_vector;
function slv_to_uint1246_t(x : std_logic_vector) return uint1246_t;
subtype int1246_t is signed(1245 downto 0);
constant int1246_t_SLV_LEN : integer := 1246;
function int1246_t_to_slv(x : int1246_t) return std_logic_vector;
function slv_to_int1246_t(x : std_logic_vector) return int1246_t;
subtype uint1247_t is unsigned(1246 downto 0);
constant uint1247_t_SLV_LEN : integer := 1247;
function uint1247_t_to_slv(x : uint1247_t) return std_logic_vector;
function slv_to_uint1247_t(x : std_logic_vector) return uint1247_t;
subtype int1247_t is signed(1246 downto 0);
constant int1247_t_SLV_LEN : integer := 1247;
function int1247_t_to_slv(x : int1247_t) return std_logic_vector;
function slv_to_int1247_t(x : std_logic_vector) return int1247_t;
subtype uint1248_t is unsigned(1247 downto 0);
constant uint1248_t_SLV_LEN : integer := 1248;
function uint1248_t_to_slv(x : uint1248_t) return std_logic_vector;
function slv_to_uint1248_t(x : std_logic_vector) return uint1248_t;
subtype int1248_t is signed(1247 downto 0);
constant int1248_t_SLV_LEN : integer := 1248;
function int1248_t_to_slv(x : int1248_t) return std_logic_vector;
function slv_to_int1248_t(x : std_logic_vector) return int1248_t;
subtype uint1249_t is unsigned(1248 downto 0);
constant uint1249_t_SLV_LEN : integer := 1249;
function uint1249_t_to_slv(x : uint1249_t) return std_logic_vector;
function slv_to_uint1249_t(x : std_logic_vector) return uint1249_t;
subtype int1249_t is signed(1248 downto 0);
constant int1249_t_SLV_LEN : integer := 1249;
function int1249_t_to_slv(x : int1249_t) return std_logic_vector;
function slv_to_int1249_t(x : std_logic_vector) return int1249_t;
subtype uint1250_t is unsigned(1249 downto 0);
constant uint1250_t_SLV_LEN : integer := 1250;
function uint1250_t_to_slv(x : uint1250_t) return std_logic_vector;
function slv_to_uint1250_t(x : std_logic_vector) return uint1250_t;
subtype int1250_t is signed(1249 downto 0);
constant int1250_t_SLV_LEN : integer := 1250;
function int1250_t_to_slv(x : int1250_t) return std_logic_vector;
function slv_to_int1250_t(x : std_logic_vector) return int1250_t;
subtype uint1251_t is unsigned(1250 downto 0);
constant uint1251_t_SLV_LEN : integer := 1251;
function uint1251_t_to_slv(x : uint1251_t) return std_logic_vector;
function slv_to_uint1251_t(x : std_logic_vector) return uint1251_t;
subtype int1251_t is signed(1250 downto 0);
constant int1251_t_SLV_LEN : integer := 1251;
function int1251_t_to_slv(x : int1251_t) return std_logic_vector;
function slv_to_int1251_t(x : std_logic_vector) return int1251_t;
subtype uint1252_t is unsigned(1251 downto 0);
constant uint1252_t_SLV_LEN : integer := 1252;
function uint1252_t_to_slv(x : uint1252_t) return std_logic_vector;
function slv_to_uint1252_t(x : std_logic_vector) return uint1252_t;
subtype int1252_t is signed(1251 downto 0);
constant int1252_t_SLV_LEN : integer := 1252;
function int1252_t_to_slv(x : int1252_t) return std_logic_vector;
function slv_to_int1252_t(x : std_logic_vector) return int1252_t;
subtype uint1253_t is unsigned(1252 downto 0);
constant uint1253_t_SLV_LEN : integer := 1253;
function uint1253_t_to_slv(x : uint1253_t) return std_logic_vector;
function slv_to_uint1253_t(x : std_logic_vector) return uint1253_t;
subtype int1253_t is signed(1252 downto 0);
constant int1253_t_SLV_LEN : integer := 1253;
function int1253_t_to_slv(x : int1253_t) return std_logic_vector;
function slv_to_int1253_t(x : std_logic_vector) return int1253_t;
subtype uint1254_t is unsigned(1253 downto 0);
constant uint1254_t_SLV_LEN : integer := 1254;
function uint1254_t_to_slv(x : uint1254_t) return std_logic_vector;
function slv_to_uint1254_t(x : std_logic_vector) return uint1254_t;
subtype int1254_t is signed(1253 downto 0);
constant int1254_t_SLV_LEN : integer := 1254;
function int1254_t_to_slv(x : int1254_t) return std_logic_vector;
function slv_to_int1254_t(x : std_logic_vector) return int1254_t;
subtype uint1255_t is unsigned(1254 downto 0);
constant uint1255_t_SLV_LEN : integer := 1255;
function uint1255_t_to_slv(x : uint1255_t) return std_logic_vector;
function slv_to_uint1255_t(x : std_logic_vector) return uint1255_t;
subtype int1255_t is signed(1254 downto 0);
constant int1255_t_SLV_LEN : integer := 1255;
function int1255_t_to_slv(x : int1255_t) return std_logic_vector;
function slv_to_int1255_t(x : std_logic_vector) return int1255_t;
subtype uint1256_t is unsigned(1255 downto 0);
constant uint1256_t_SLV_LEN : integer := 1256;
function uint1256_t_to_slv(x : uint1256_t) return std_logic_vector;
function slv_to_uint1256_t(x : std_logic_vector) return uint1256_t;
subtype int1256_t is signed(1255 downto 0);
constant int1256_t_SLV_LEN : integer := 1256;
function int1256_t_to_slv(x : int1256_t) return std_logic_vector;
function slv_to_int1256_t(x : std_logic_vector) return int1256_t;
subtype uint1257_t is unsigned(1256 downto 0);
constant uint1257_t_SLV_LEN : integer := 1257;
function uint1257_t_to_slv(x : uint1257_t) return std_logic_vector;
function slv_to_uint1257_t(x : std_logic_vector) return uint1257_t;
subtype int1257_t is signed(1256 downto 0);
constant int1257_t_SLV_LEN : integer := 1257;
function int1257_t_to_slv(x : int1257_t) return std_logic_vector;
function slv_to_int1257_t(x : std_logic_vector) return int1257_t;
subtype uint1258_t is unsigned(1257 downto 0);
constant uint1258_t_SLV_LEN : integer := 1258;
function uint1258_t_to_slv(x : uint1258_t) return std_logic_vector;
function slv_to_uint1258_t(x : std_logic_vector) return uint1258_t;
subtype int1258_t is signed(1257 downto 0);
constant int1258_t_SLV_LEN : integer := 1258;
function int1258_t_to_slv(x : int1258_t) return std_logic_vector;
function slv_to_int1258_t(x : std_logic_vector) return int1258_t;
subtype uint1259_t is unsigned(1258 downto 0);
constant uint1259_t_SLV_LEN : integer := 1259;
function uint1259_t_to_slv(x : uint1259_t) return std_logic_vector;
function slv_to_uint1259_t(x : std_logic_vector) return uint1259_t;
subtype int1259_t is signed(1258 downto 0);
constant int1259_t_SLV_LEN : integer := 1259;
function int1259_t_to_slv(x : int1259_t) return std_logic_vector;
function slv_to_int1259_t(x : std_logic_vector) return int1259_t;
subtype uint1260_t is unsigned(1259 downto 0);
constant uint1260_t_SLV_LEN : integer := 1260;
function uint1260_t_to_slv(x : uint1260_t) return std_logic_vector;
function slv_to_uint1260_t(x : std_logic_vector) return uint1260_t;
subtype int1260_t is signed(1259 downto 0);
constant int1260_t_SLV_LEN : integer := 1260;
function int1260_t_to_slv(x : int1260_t) return std_logic_vector;
function slv_to_int1260_t(x : std_logic_vector) return int1260_t;
subtype uint1261_t is unsigned(1260 downto 0);
constant uint1261_t_SLV_LEN : integer := 1261;
function uint1261_t_to_slv(x : uint1261_t) return std_logic_vector;
function slv_to_uint1261_t(x : std_logic_vector) return uint1261_t;
subtype int1261_t is signed(1260 downto 0);
constant int1261_t_SLV_LEN : integer := 1261;
function int1261_t_to_slv(x : int1261_t) return std_logic_vector;
function slv_to_int1261_t(x : std_logic_vector) return int1261_t;
subtype uint1262_t is unsigned(1261 downto 0);
constant uint1262_t_SLV_LEN : integer := 1262;
function uint1262_t_to_slv(x : uint1262_t) return std_logic_vector;
function slv_to_uint1262_t(x : std_logic_vector) return uint1262_t;
subtype int1262_t is signed(1261 downto 0);
constant int1262_t_SLV_LEN : integer := 1262;
function int1262_t_to_slv(x : int1262_t) return std_logic_vector;
function slv_to_int1262_t(x : std_logic_vector) return int1262_t;
subtype uint1263_t is unsigned(1262 downto 0);
constant uint1263_t_SLV_LEN : integer := 1263;
function uint1263_t_to_slv(x : uint1263_t) return std_logic_vector;
function slv_to_uint1263_t(x : std_logic_vector) return uint1263_t;
subtype int1263_t is signed(1262 downto 0);
constant int1263_t_SLV_LEN : integer := 1263;
function int1263_t_to_slv(x : int1263_t) return std_logic_vector;
function slv_to_int1263_t(x : std_logic_vector) return int1263_t;
subtype uint1264_t is unsigned(1263 downto 0);
constant uint1264_t_SLV_LEN : integer := 1264;
function uint1264_t_to_slv(x : uint1264_t) return std_logic_vector;
function slv_to_uint1264_t(x : std_logic_vector) return uint1264_t;
subtype int1264_t is signed(1263 downto 0);
constant int1264_t_SLV_LEN : integer := 1264;
function int1264_t_to_slv(x : int1264_t) return std_logic_vector;
function slv_to_int1264_t(x : std_logic_vector) return int1264_t;
subtype uint1265_t is unsigned(1264 downto 0);
constant uint1265_t_SLV_LEN : integer := 1265;
function uint1265_t_to_slv(x : uint1265_t) return std_logic_vector;
function slv_to_uint1265_t(x : std_logic_vector) return uint1265_t;
subtype int1265_t is signed(1264 downto 0);
constant int1265_t_SLV_LEN : integer := 1265;
function int1265_t_to_slv(x : int1265_t) return std_logic_vector;
function slv_to_int1265_t(x : std_logic_vector) return int1265_t;
subtype uint1266_t is unsigned(1265 downto 0);
constant uint1266_t_SLV_LEN : integer := 1266;
function uint1266_t_to_slv(x : uint1266_t) return std_logic_vector;
function slv_to_uint1266_t(x : std_logic_vector) return uint1266_t;
subtype int1266_t is signed(1265 downto 0);
constant int1266_t_SLV_LEN : integer := 1266;
function int1266_t_to_slv(x : int1266_t) return std_logic_vector;
function slv_to_int1266_t(x : std_logic_vector) return int1266_t;
subtype uint1267_t is unsigned(1266 downto 0);
constant uint1267_t_SLV_LEN : integer := 1267;
function uint1267_t_to_slv(x : uint1267_t) return std_logic_vector;
function slv_to_uint1267_t(x : std_logic_vector) return uint1267_t;
subtype int1267_t is signed(1266 downto 0);
constant int1267_t_SLV_LEN : integer := 1267;
function int1267_t_to_slv(x : int1267_t) return std_logic_vector;
function slv_to_int1267_t(x : std_logic_vector) return int1267_t;
subtype uint1268_t is unsigned(1267 downto 0);
constant uint1268_t_SLV_LEN : integer := 1268;
function uint1268_t_to_slv(x : uint1268_t) return std_logic_vector;
function slv_to_uint1268_t(x : std_logic_vector) return uint1268_t;
subtype int1268_t is signed(1267 downto 0);
constant int1268_t_SLV_LEN : integer := 1268;
function int1268_t_to_slv(x : int1268_t) return std_logic_vector;
function slv_to_int1268_t(x : std_logic_vector) return int1268_t;
subtype uint1269_t is unsigned(1268 downto 0);
constant uint1269_t_SLV_LEN : integer := 1269;
function uint1269_t_to_slv(x : uint1269_t) return std_logic_vector;
function slv_to_uint1269_t(x : std_logic_vector) return uint1269_t;
subtype int1269_t is signed(1268 downto 0);
constant int1269_t_SLV_LEN : integer := 1269;
function int1269_t_to_slv(x : int1269_t) return std_logic_vector;
function slv_to_int1269_t(x : std_logic_vector) return int1269_t;
subtype uint1270_t is unsigned(1269 downto 0);
constant uint1270_t_SLV_LEN : integer := 1270;
function uint1270_t_to_slv(x : uint1270_t) return std_logic_vector;
function slv_to_uint1270_t(x : std_logic_vector) return uint1270_t;
subtype int1270_t is signed(1269 downto 0);
constant int1270_t_SLV_LEN : integer := 1270;
function int1270_t_to_slv(x : int1270_t) return std_logic_vector;
function slv_to_int1270_t(x : std_logic_vector) return int1270_t;
subtype uint1271_t is unsigned(1270 downto 0);
constant uint1271_t_SLV_LEN : integer := 1271;
function uint1271_t_to_slv(x : uint1271_t) return std_logic_vector;
function slv_to_uint1271_t(x : std_logic_vector) return uint1271_t;
subtype int1271_t is signed(1270 downto 0);
constant int1271_t_SLV_LEN : integer := 1271;
function int1271_t_to_slv(x : int1271_t) return std_logic_vector;
function slv_to_int1271_t(x : std_logic_vector) return int1271_t;
subtype uint1272_t is unsigned(1271 downto 0);
constant uint1272_t_SLV_LEN : integer := 1272;
function uint1272_t_to_slv(x : uint1272_t) return std_logic_vector;
function slv_to_uint1272_t(x : std_logic_vector) return uint1272_t;
subtype int1272_t is signed(1271 downto 0);
constant int1272_t_SLV_LEN : integer := 1272;
function int1272_t_to_slv(x : int1272_t) return std_logic_vector;
function slv_to_int1272_t(x : std_logic_vector) return int1272_t;
subtype uint1273_t is unsigned(1272 downto 0);
constant uint1273_t_SLV_LEN : integer := 1273;
function uint1273_t_to_slv(x : uint1273_t) return std_logic_vector;
function slv_to_uint1273_t(x : std_logic_vector) return uint1273_t;
subtype int1273_t is signed(1272 downto 0);
constant int1273_t_SLV_LEN : integer := 1273;
function int1273_t_to_slv(x : int1273_t) return std_logic_vector;
function slv_to_int1273_t(x : std_logic_vector) return int1273_t;
subtype uint1274_t is unsigned(1273 downto 0);
constant uint1274_t_SLV_LEN : integer := 1274;
function uint1274_t_to_slv(x : uint1274_t) return std_logic_vector;
function slv_to_uint1274_t(x : std_logic_vector) return uint1274_t;
subtype int1274_t is signed(1273 downto 0);
constant int1274_t_SLV_LEN : integer := 1274;
function int1274_t_to_slv(x : int1274_t) return std_logic_vector;
function slv_to_int1274_t(x : std_logic_vector) return int1274_t;
subtype uint1275_t is unsigned(1274 downto 0);
constant uint1275_t_SLV_LEN : integer := 1275;
function uint1275_t_to_slv(x : uint1275_t) return std_logic_vector;
function slv_to_uint1275_t(x : std_logic_vector) return uint1275_t;
subtype int1275_t is signed(1274 downto 0);
constant int1275_t_SLV_LEN : integer := 1275;
function int1275_t_to_slv(x : int1275_t) return std_logic_vector;
function slv_to_int1275_t(x : std_logic_vector) return int1275_t;
subtype uint1276_t is unsigned(1275 downto 0);
constant uint1276_t_SLV_LEN : integer := 1276;
function uint1276_t_to_slv(x : uint1276_t) return std_logic_vector;
function slv_to_uint1276_t(x : std_logic_vector) return uint1276_t;
subtype int1276_t is signed(1275 downto 0);
constant int1276_t_SLV_LEN : integer := 1276;
function int1276_t_to_slv(x : int1276_t) return std_logic_vector;
function slv_to_int1276_t(x : std_logic_vector) return int1276_t;
subtype uint1277_t is unsigned(1276 downto 0);
constant uint1277_t_SLV_LEN : integer := 1277;
function uint1277_t_to_slv(x : uint1277_t) return std_logic_vector;
function slv_to_uint1277_t(x : std_logic_vector) return uint1277_t;
subtype int1277_t is signed(1276 downto 0);
constant int1277_t_SLV_LEN : integer := 1277;
function int1277_t_to_slv(x : int1277_t) return std_logic_vector;
function slv_to_int1277_t(x : std_logic_vector) return int1277_t;
subtype uint1278_t is unsigned(1277 downto 0);
constant uint1278_t_SLV_LEN : integer := 1278;
function uint1278_t_to_slv(x : uint1278_t) return std_logic_vector;
function slv_to_uint1278_t(x : std_logic_vector) return uint1278_t;
subtype int1278_t is signed(1277 downto 0);
constant int1278_t_SLV_LEN : integer := 1278;
function int1278_t_to_slv(x : int1278_t) return std_logic_vector;
function slv_to_int1278_t(x : std_logic_vector) return int1278_t;
subtype uint1279_t is unsigned(1278 downto 0);
constant uint1279_t_SLV_LEN : integer := 1279;
function uint1279_t_to_slv(x : uint1279_t) return std_logic_vector;
function slv_to_uint1279_t(x : std_logic_vector) return uint1279_t;
subtype int1279_t is signed(1278 downto 0);
constant int1279_t_SLV_LEN : integer := 1279;
function int1279_t_to_slv(x : int1279_t) return std_logic_vector;
function slv_to_int1279_t(x : std_logic_vector) return int1279_t;
subtype uint1280_t is unsigned(1279 downto 0);
constant uint1280_t_SLV_LEN : integer := 1280;
function uint1280_t_to_slv(x : uint1280_t) return std_logic_vector;
function slv_to_uint1280_t(x : std_logic_vector) return uint1280_t;
subtype int1280_t is signed(1279 downto 0);
constant int1280_t_SLV_LEN : integer := 1280;
function int1280_t_to_slv(x : int1280_t) return std_logic_vector;
function slv_to_int1280_t(x : std_logic_vector) return int1280_t;
subtype uint1281_t is unsigned(1280 downto 0);
constant uint1281_t_SLV_LEN : integer := 1281;
function uint1281_t_to_slv(x : uint1281_t) return std_logic_vector;
function slv_to_uint1281_t(x : std_logic_vector) return uint1281_t;
subtype int1281_t is signed(1280 downto 0);
constant int1281_t_SLV_LEN : integer := 1281;
function int1281_t_to_slv(x : int1281_t) return std_logic_vector;
function slv_to_int1281_t(x : std_logic_vector) return int1281_t;
subtype uint1282_t is unsigned(1281 downto 0);
constant uint1282_t_SLV_LEN : integer := 1282;
function uint1282_t_to_slv(x : uint1282_t) return std_logic_vector;
function slv_to_uint1282_t(x : std_logic_vector) return uint1282_t;
subtype int1282_t is signed(1281 downto 0);
constant int1282_t_SLV_LEN : integer := 1282;
function int1282_t_to_slv(x : int1282_t) return std_logic_vector;
function slv_to_int1282_t(x : std_logic_vector) return int1282_t;
subtype uint1283_t is unsigned(1282 downto 0);
constant uint1283_t_SLV_LEN : integer := 1283;
function uint1283_t_to_slv(x : uint1283_t) return std_logic_vector;
function slv_to_uint1283_t(x : std_logic_vector) return uint1283_t;
subtype int1283_t is signed(1282 downto 0);
constant int1283_t_SLV_LEN : integer := 1283;
function int1283_t_to_slv(x : int1283_t) return std_logic_vector;
function slv_to_int1283_t(x : std_logic_vector) return int1283_t;
subtype uint1284_t is unsigned(1283 downto 0);
constant uint1284_t_SLV_LEN : integer := 1284;
function uint1284_t_to_slv(x : uint1284_t) return std_logic_vector;
function slv_to_uint1284_t(x : std_logic_vector) return uint1284_t;
subtype int1284_t is signed(1283 downto 0);
constant int1284_t_SLV_LEN : integer := 1284;
function int1284_t_to_slv(x : int1284_t) return std_logic_vector;
function slv_to_int1284_t(x : std_logic_vector) return int1284_t;
subtype uint1285_t is unsigned(1284 downto 0);
constant uint1285_t_SLV_LEN : integer := 1285;
function uint1285_t_to_slv(x : uint1285_t) return std_logic_vector;
function slv_to_uint1285_t(x : std_logic_vector) return uint1285_t;
subtype int1285_t is signed(1284 downto 0);
constant int1285_t_SLV_LEN : integer := 1285;
function int1285_t_to_slv(x : int1285_t) return std_logic_vector;
function slv_to_int1285_t(x : std_logic_vector) return int1285_t;
subtype uint1286_t is unsigned(1285 downto 0);
constant uint1286_t_SLV_LEN : integer := 1286;
function uint1286_t_to_slv(x : uint1286_t) return std_logic_vector;
function slv_to_uint1286_t(x : std_logic_vector) return uint1286_t;
subtype int1286_t is signed(1285 downto 0);
constant int1286_t_SLV_LEN : integer := 1286;
function int1286_t_to_slv(x : int1286_t) return std_logic_vector;
function slv_to_int1286_t(x : std_logic_vector) return int1286_t;
subtype uint1287_t is unsigned(1286 downto 0);
constant uint1287_t_SLV_LEN : integer := 1287;
function uint1287_t_to_slv(x : uint1287_t) return std_logic_vector;
function slv_to_uint1287_t(x : std_logic_vector) return uint1287_t;
subtype int1287_t is signed(1286 downto 0);
constant int1287_t_SLV_LEN : integer := 1287;
function int1287_t_to_slv(x : int1287_t) return std_logic_vector;
function slv_to_int1287_t(x : std_logic_vector) return int1287_t;
subtype uint1288_t is unsigned(1287 downto 0);
constant uint1288_t_SLV_LEN : integer := 1288;
function uint1288_t_to_slv(x : uint1288_t) return std_logic_vector;
function slv_to_uint1288_t(x : std_logic_vector) return uint1288_t;
subtype int1288_t is signed(1287 downto 0);
constant int1288_t_SLV_LEN : integer := 1288;
function int1288_t_to_slv(x : int1288_t) return std_logic_vector;
function slv_to_int1288_t(x : std_logic_vector) return int1288_t;
subtype uint1289_t is unsigned(1288 downto 0);
constant uint1289_t_SLV_LEN : integer := 1289;
function uint1289_t_to_slv(x : uint1289_t) return std_logic_vector;
function slv_to_uint1289_t(x : std_logic_vector) return uint1289_t;
subtype int1289_t is signed(1288 downto 0);
constant int1289_t_SLV_LEN : integer := 1289;
function int1289_t_to_slv(x : int1289_t) return std_logic_vector;
function slv_to_int1289_t(x : std_logic_vector) return int1289_t;
subtype uint1290_t is unsigned(1289 downto 0);
constant uint1290_t_SLV_LEN : integer := 1290;
function uint1290_t_to_slv(x : uint1290_t) return std_logic_vector;
function slv_to_uint1290_t(x : std_logic_vector) return uint1290_t;
subtype int1290_t is signed(1289 downto 0);
constant int1290_t_SLV_LEN : integer := 1290;
function int1290_t_to_slv(x : int1290_t) return std_logic_vector;
function slv_to_int1290_t(x : std_logic_vector) return int1290_t;
subtype uint1291_t is unsigned(1290 downto 0);
constant uint1291_t_SLV_LEN : integer := 1291;
function uint1291_t_to_slv(x : uint1291_t) return std_logic_vector;
function slv_to_uint1291_t(x : std_logic_vector) return uint1291_t;
subtype int1291_t is signed(1290 downto 0);
constant int1291_t_SLV_LEN : integer := 1291;
function int1291_t_to_slv(x : int1291_t) return std_logic_vector;
function slv_to_int1291_t(x : std_logic_vector) return int1291_t;
subtype uint1292_t is unsigned(1291 downto 0);
constant uint1292_t_SLV_LEN : integer := 1292;
function uint1292_t_to_slv(x : uint1292_t) return std_logic_vector;
function slv_to_uint1292_t(x : std_logic_vector) return uint1292_t;
subtype int1292_t is signed(1291 downto 0);
constant int1292_t_SLV_LEN : integer := 1292;
function int1292_t_to_slv(x : int1292_t) return std_logic_vector;
function slv_to_int1292_t(x : std_logic_vector) return int1292_t;
subtype uint1293_t is unsigned(1292 downto 0);
constant uint1293_t_SLV_LEN : integer := 1293;
function uint1293_t_to_slv(x : uint1293_t) return std_logic_vector;
function slv_to_uint1293_t(x : std_logic_vector) return uint1293_t;
subtype int1293_t is signed(1292 downto 0);
constant int1293_t_SLV_LEN : integer := 1293;
function int1293_t_to_slv(x : int1293_t) return std_logic_vector;
function slv_to_int1293_t(x : std_logic_vector) return int1293_t;
subtype uint1294_t is unsigned(1293 downto 0);
constant uint1294_t_SLV_LEN : integer := 1294;
function uint1294_t_to_slv(x : uint1294_t) return std_logic_vector;
function slv_to_uint1294_t(x : std_logic_vector) return uint1294_t;
subtype int1294_t is signed(1293 downto 0);
constant int1294_t_SLV_LEN : integer := 1294;
function int1294_t_to_slv(x : int1294_t) return std_logic_vector;
function slv_to_int1294_t(x : std_logic_vector) return int1294_t;
subtype uint1295_t is unsigned(1294 downto 0);
constant uint1295_t_SLV_LEN : integer := 1295;
function uint1295_t_to_slv(x : uint1295_t) return std_logic_vector;
function slv_to_uint1295_t(x : std_logic_vector) return uint1295_t;
subtype int1295_t is signed(1294 downto 0);
constant int1295_t_SLV_LEN : integer := 1295;
function int1295_t_to_slv(x : int1295_t) return std_logic_vector;
function slv_to_int1295_t(x : std_logic_vector) return int1295_t;
subtype uint1296_t is unsigned(1295 downto 0);
constant uint1296_t_SLV_LEN : integer := 1296;
function uint1296_t_to_slv(x : uint1296_t) return std_logic_vector;
function slv_to_uint1296_t(x : std_logic_vector) return uint1296_t;
subtype int1296_t is signed(1295 downto 0);
constant int1296_t_SLV_LEN : integer := 1296;
function int1296_t_to_slv(x : int1296_t) return std_logic_vector;
function slv_to_int1296_t(x : std_logic_vector) return int1296_t;
subtype uint1297_t is unsigned(1296 downto 0);
constant uint1297_t_SLV_LEN : integer := 1297;
function uint1297_t_to_slv(x : uint1297_t) return std_logic_vector;
function slv_to_uint1297_t(x : std_logic_vector) return uint1297_t;
subtype int1297_t is signed(1296 downto 0);
constant int1297_t_SLV_LEN : integer := 1297;
function int1297_t_to_slv(x : int1297_t) return std_logic_vector;
function slv_to_int1297_t(x : std_logic_vector) return int1297_t;
subtype uint1298_t is unsigned(1297 downto 0);
constant uint1298_t_SLV_LEN : integer := 1298;
function uint1298_t_to_slv(x : uint1298_t) return std_logic_vector;
function slv_to_uint1298_t(x : std_logic_vector) return uint1298_t;
subtype int1298_t is signed(1297 downto 0);
constant int1298_t_SLV_LEN : integer := 1298;
function int1298_t_to_slv(x : int1298_t) return std_logic_vector;
function slv_to_int1298_t(x : std_logic_vector) return int1298_t;
subtype uint1299_t is unsigned(1298 downto 0);
constant uint1299_t_SLV_LEN : integer := 1299;
function uint1299_t_to_slv(x : uint1299_t) return std_logic_vector;
function slv_to_uint1299_t(x : std_logic_vector) return uint1299_t;
subtype int1299_t is signed(1298 downto 0);
constant int1299_t_SLV_LEN : integer := 1299;
function int1299_t_to_slv(x : int1299_t) return std_logic_vector;
function slv_to_int1299_t(x : std_logic_vector) return int1299_t;
subtype uint1300_t is unsigned(1299 downto 0);
constant uint1300_t_SLV_LEN : integer := 1300;
function uint1300_t_to_slv(x : uint1300_t) return std_logic_vector;
function slv_to_uint1300_t(x : std_logic_vector) return uint1300_t;
subtype int1300_t is signed(1299 downto 0);
constant int1300_t_SLV_LEN : integer := 1300;
function int1300_t_to_slv(x : int1300_t) return std_logic_vector;
function slv_to_int1300_t(x : std_logic_vector) return int1300_t;
subtype uint1301_t is unsigned(1300 downto 0);
constant uint1301_t_SLV_LEN : integer := 1301;
function uint1301_t_to_slv(x : uint1301_t) return std_logic_vector;
function slv_to_uint1301_t(x : std_logic_vector) return uint1301_t;
subtype int1301_t is signed(1300 downto 0);
constant int1301_t_SLV_LEN : integer := 1301;
function int1301_t_to_slv(x : int1301_t) return std_logic_vector;
function slv_to_int1301_t(x : std_logic_vector) return int1301_t;
subtype uint1302_t is unsigned(1301 downto 0);
constant uint1302_t_SLV_LEN : integer := 1302;
function uint1302_t_to_slv(x : uint1302_t) return std_logic_vector;
function slv_to_uint1302_t(x : std_logic_vector) return uint1302_t;
subtype int1302_t is signed(1301 downto 0);
constant int1302_t_SLV_LEN : integer := 1302;
function int1302_t_to_slv(x : int1302_t) return std_logic_vector;
function slv_to_int1302_t(x : std_logic_vector) return int1302_t;
subtype uint1303_t is unsigned(1302 downto 0);
constant uint1303_t_SLV_LEN : integer := 1303;
function uint1303_t_to_slv(x : uint1303_t) return std_logic_vector;
function slv_to_uint1303_t(x : std_logic_vector) return uint1303_t;
subtype int1303_t is signed(1302 downto 0);
constant int1303_t_SLV_LEN : integer := 1303;
function int1303_t_to_slv(x : int1303_t) return std_logic_vector;
function slv_to_int1303_t(x : std_logic_vector) return int1303_t;
subtype uint1304_t is unsigned(1303 downto 0);
constant uint1304_t_SLV_LEN : integer := 1304;
function uint1304_t_to_slv(x : uint1304_t) return std_logic_vector;
function slv_to_uint1304_t(x : std_logic_vector) return uint1304_t;
subtype int1304_t is signed(1303 downto 0);
constant int1304_t_SLV_LEN : integer := 1304;
function int1304_t_to_slv(x : int1304_t) return std_logic_vector;
function slv_to_int1304_t(x : std_logic_vector) return int1304_t;
subtype uint1305_t is unsigned(1304 downto 0);
constant uint1305_t_SLV_LEN : integer := 1305;
function uint1305_t_to_slv(x : uint1305_t) return std_logic_vector;
function slv_to_uint1305_t(x : std_logic_vector) return uint1305_t;
subtype int1305_t is signed(1304 downto 0);
constant int1305_t_SLV_LEN : integer := 1305;
function int1305_t_to_slv(x : int1305_t) return std_logic_vector;
function slv_to_int1305_t(x : std_logic_vector) return int1305_t;
subtype uint1306_t is unsigned(1305 downto 0);
constant uint1306_t_SLV_LEN : integer := 1306;
function uint1306_t_to_slv(x : uint1306_t) return std_logic_vector;
function slv_to_uint1306_t(x : std_logic_vector) return uint1306_t;
subtype int1306_t is signed(1305 downto 0);
constant int1306_t_SLV_LEN : integer := 1306;
function int1306_t_to_slv(x : int1306_t) return std_logic_vector;
function slv_to_int1306_t(x : std_logic_vector) return int1306_t;
subtype uint1307_t is unsigned(1306 downto 0);
constant uint1307_t_SLV_LEN : integer := 1307;
function uint1307_t_to_slv(x : uint1307_t) return std_logic_vector;
function slv_to_uint1307_t(x : std_logic_vector) return uint1307_t;
subtype int1307_t is signed(1306 downto 0);
constant int1307_t_SLV_LEN : integer := 1307;
function int1307_t_to_slv(x : int1307_t) return std_logic_vector;
function slv_to_int1307_t(x : std_logic_vector) return int1307_t;
subtype uint1308_t is unsigned(1307 downto 0);
constant uint1308_t_SLV_LEN : integer := 1308;
function uint1308_t_to_slv(x : uint1308_t) return std_logic_vector;
function slv_to_uint1308_t(x : std_logic_vector) return uint1308_t;
subtype int1308_t is signed(1307 downto 0);
constant int1308_t_SLV_LEN : integer := 1308;
function int1308_t_to_slv(x : int1308_t) return std_logic_vector;
function slv_to_int1308_t(x : std_logic_vector) return int1308_t;
subtype uint1309_t is unsigned(1308 downto 0);
constant uint1309_t_SLV_LEN : integer := 1309;
function uint1309_t_to_slv(x : uint1309_t) return std_logic_vector;
function slv_to_uint1309_t(x : std_logic_vector) return uint1309_t;
subtype int1309_t is signed(1308 downto 0);
constant int1309_t_SLV_LEN : integer := 1309;
function int1309_t_to_slv(x : int1309_t) return std_logic_vector;
function slv_to_int1309_t(x : std_logic_vector) return int1309_t;
subtype uint1310_t is unsigned(1309 downto 0);
constant uint1310_t_SLV_LEN : integer := 1310;
function uint1310_t_to_slv(x : uint1310_t) return std_logic_vector;
function slv_to_uint1310_t(x : std_logic_vector) return uint1310_t;
subtype int1310_t is signed(1309 downto 0);
constant int1310_t_SLV_LEN : integer := 1310;
function int1310_t_to_slv(x : int1310_t) return std_logic_vector;
function slv_to_int1310_t(x : std_logic_vector) return int1310_t;
subtype uint1311_t is unsigned(1310 downto 0);
constant uint1311_t_SLV_LEN : integer := 1311;
function uint1311_t_to_slv(x : uint1311_t) return std_logic_vector;
function slv_to_uint1311_t(x : std_logic_vector) return uint1311_t;
subtype int1311_t is signed(1310 downto 0);
constant int1311_t_SLV_LEN : integer := 1311;
function int1311_t_to_slv(x : int1311_t) return std_logic_vector;
function slv_to_int1311_t(x : std_logic_vector) return int1311_t;
subtype uint1312_t is unsigned(1311 downto 0);
constant uint1312_t_SLV_LEN : integer := 1312;
function uint1312_t_to_slv(x : uint1312_t) return std_logic_vector;
function slv_to_uint1312_t(x : std_logic_vector) return uint1312_t;
subtype int1312_t is signed(1311 downto 0);
constant int1312_t_SLV_LEN : integer := 1312;
function int1312_t_to_slv(x : int1312_t) return std_logic_vector;
function slv_to_int1312_t(x : std_logic_vector) return int1312_t;
subtype uint1313_t is unsigned(1312 downto 0);
constant uint1313_t_SLV_LEN : integer := 1313;
function uint1313_t_to_slv(x : uint1313_t) return std_logic_vector;
function slv_to_uint1313_t(x : std_logic_vector) return uint1313_t;
subtype int1313_t is signed(1312 downto 0);
constant int1313_t_SLV_LEN : integer := 1313;
function int1313_t_to_slv(x : int1313_t) return std_logic_vector;
function slv_to_int1313_t(x : std_logic_vector) return int1313_t;
subtype uint1314_t is unsigned(1313 downto 0);
constant uint1314_t_SLV_LEN : integer := 1314;
function uint1314_t_to_slv(x : uint1314_t) return std_logic_vector;
function slv_to_uint1314_t(x : std_logic_vector) return uint1314_t;
subtype int1314_t is signed(1313 downto 0);
constant int1314_t_SLV_LEN : integer := 1314;
function int1314_t_to_slv(x : int1314_t) return std_logic_vector;
function slv_to_int1314_t(x : std_logic_vector) return int1314_t;
subtype uint1315_t is unsigned(1314 downto 0);
constant uint1315_t_SLV_LEN : integer := 1315;
function uint1315_t_to_slv(x : uint1315_t) return std_logic_vector;
function slv_to_uint1315_t(x : std_logic_vector) return uint1315_t;
subtype int1315_t is signed(1314 downto 0);
constant int1315_t_SLV_LEN : integer := 1315;
function int1315_t_to_slv(x : int1315_t) return std_logic_vector;
function slv_to_int1315_t(x : std_logic_vector) return int1315_t;
subtype uint1316_t is unsigned(1315 downto 0);
constant uint1316_t_SLV_LEN : integer := 1316;
function uint1316_t_to_slv(x : uint1316_t) return std_logic_vector;
function slv_to_uint1316_t(x : std_logic_vector) return uint1316_t;
subtype int1316_t is signed(1315 downto 0);
constant int1316_t_SLV_LEN : integer := 1316;
function int1316_t_to_slv(x : int1316_t) return std_logic_vector;
function slv_to_int1316_t(x : std_logic_vector) return int1316_t;
subtype uint1317_t is unsigned(1316 downto 0);
constant uint1317_t_SLV_LEN : integer := 1317;
function uint1317_t_to_slv(x : uint1317_t) return std_logic_vector;
function slv_to_uint1317_t(x : std_logic_vector) return uint1317_t;
subtype int1317_t is signed(1316 downto 0);
constant int1317_t_SLV_LEN : integer := 1317;
function int1317_t_to_slv(x : int1317_t) return std_logic_vector;
function slv_to_int1317_t(x : std_logic_vector) return int1317_t;
subtype uint1318_t is unsigned(1317 downto 0);
constant uint1318_t_SLV_LEN : integer := 1318;
function uint1318_t_to_slv(x : uint1318_t) return std_logic_vector;
function slv_to_uint1318_t(x : std_logic_vector) return uint1318_t;
subtype int1318_t is signed(1317 downto 0);
constant int1318_t_SLV_LEN : integer := 1318;
function int1318_t_to_slv(x : int1318_t) return std_logic_vector;
function slv_to_int1318_t(x : std_logic_vector) return int1318_t;
subtype uint1319_t is unsigned(1318 downto 0);
constant uint1319_t_SLV_LEN : integer := 1319;
function uint1319_t_to_slv(x : uint1319_t) return std_logic_vector;
function slv_to_uint1319_t(x : std_logic_vector) return uint1319_t;
subtype int1319_t is signed(1318 downto 0);
constant int1319_t_SLV_LEN : integer := 1319;
function int1319_t_to_slv(x : int1319_t) return std_logic_vector;
function slv_to_int1319_t(x : std_logic_vector) return int1319_t;
subtype uint1320_t is unsigned(1319 downto 0);
constant uint1320_t_SLV_LEN : integer := 1320;
function uint1320_t_to_slv(x : uint1320_t) return std_logic_vector;
function slv_to_uint1320_t(x : std_logic_vector) return uint1320_t;
subtype int1320_t is signed(1319 downto 0);
constant int1320_t_SLV_LEN : integer := 1320;
function int1320_t_to_slv(x : int1320_t) return std_logic_vector;
function slv_to_int1320_t(x : std_logic_vector) return int1320_t;
subtype uint1321_t is unsigned(1320 downto 0);
constant uint1321_t_SLV_LEN : integer := 1321;
function uint1321_t_to_slv(x : uint1321_t) return std_logic_vector;
function slv_to_uint1321_t(x : std_logic_vector) return uint1321_t;
subtype int1321_t is signed(1320 downto 0);
constant int1321_t_SLV_LEN : integer := 1321;
function int1321_t_to_slv(x : int1321_t) return std_logic_vector;
function slv_to_int1321_t(x : std_logic_vector) return int1321_t;
subtype uint1322_t is unsigned(1321 downto 0);
constant uint1322_t_SLV_LEN : integer := 1322;
function uint1322_t_to_slv(x : uint1322_t) return std_logic_vector;
function slv_to_uint1322_t(x : std_logic_vector) return uint1322_t;
subtype int1322_t is signed(1321 downto 0);
constant int1322_t_SLV_LEN : integer := 1322;
function int1322_t_to_slv(x : int1322_t) return std_logic_vector;
function slv_to_int1322_t(x : std_logic_vector) return int1322_t;
subtype uint1323_t is unsigned(1322 downto 0);
constant uint1323_t_SLV_LEN : integer := 1323;
function uint1323_t_to_slv(x : uint1323_t) return std_logic_vector;
function slv_to_uint1323_t(x : std_logic_vector) return uint1323_t;
subtype int1323_t is signed(1322 downto 0);
constant int1323_t_SLV_LEN : integer := 1323;
function int1323_t_to_slv(x : int1323_t) return std_logic_vector;
function slv_to_int1323_t(x : std_logic_vector) return int1323_t;
subtype uint1324_t is unsigned(1323 downto 0);
constant uint1324_t_SLV_LEN : integer := 1324;
function uint1324_t_to_slv(x : uint1324_t) return std_logic_vector;
function slv_to_uint1324_t(x : std_logic_vector) return uint1324_t;
subtype int1324_t is signed(1323 downto 0);
constant int1324_t_SLV_LEN : integer := 1324;
function int1324_t_to_slv(x : int1324_t) return std_logic_vector;
function slv_to_int1324_t(x : std_logic_vector) return int1324_t;
subtype uint1325_t is unsigned(1324 downto 0);
constant uint1325_t_SLV_LEN : integer := 1325;
function uint1325_t_to_slv(x : uint1325_t) return std_logic_vector;
function slv_to_uint1325_t(x : std_logic_vector) return uint1325_t;
subtype int1325_t is signed(1324 downto 0);
constant int1325_t_SLV_LEN : integer := 1325;
function int1325_t_to_slv(x : int1325_t) return std_logic_vector;
function slv_to_int1325_t(x : std_logic_vector) return int1325_t;
subtype uint1326_t is unsigned(1325 downto 0);
constant uint1326_t_SLV_LEN : integer := 1326;
function uint1326_t_to_slv(x : uint1326_t) return std_logic_vector;
function slv_to_uint1326_t(x : std_logic_vector) return uint1326_t;
subtype int1326_t is signed(1325 downto 0);
constant int1326_t_SLV_LEN : integer := 1326;
function int1326_t_to_slv(x : int1326_t) return std_logic_vector;
function slv_to_int1326_t(x : std_logic_vector) return int1326_t;
subtype uint1327_t is unsigned(1326 downto 0);
constant uint1327_t_SLV_LEN : integer := 1327;
function uint1327_t_to_slv(x : uint1327_t) return std_logic_vector;
function slv_to_uint1327_t(x : std_logic_vector) return uint1327_t;
subtype int1327_t is signed(1326 downto 0);
constant int1327_t_SLV_LEN : integer := 1327;
function int1327_t_to_slv(x : int1327_t) return std_logic_vector;
function slv_to_int1327_t(x : std_logic_vector) return int1327_t;
subtype uint1328_t is unsigned(1327 downto 0);
constant uint1328_t_SLV_LEN : integer := 1328;
function uint1328_t_to_slv(x : uint1328_t) return std_logic_vector;
function slv_to_uint1328_t(x : std_logic_vector) return uint1328_t;
subtype int1328_t is signed(1327 downto 0);
constant int1328_t_SLV_LEN : integer := 1328;
function int1328_t_to_slv(x : int1328_t) return std_logic_vector;
function slv_to_int1328_t(x : std_logic_vector) return int1328_t;
subtype uint1329_t is unsigned(1328 downto 0);
constant uint1329_t_SLV_LEN : integer := 1329;
function uint1329_t_to_slv(x : uint1329_t) return std_logic_vector;
function slv_to_uint1329_t(x : std_logic_vector) return uint1329_t;
subtype int1329_t is signed(1328 downto 0);
constant int1329_t_SLV_LEN : integer := 1329;
function int1329_t_to_slv(x : int1329_t) return std_logic_vector;
function slv_to_int1329_t(x : std_logic_vector) return int1329_t;
subtype uint1330_t is unsigned(1329 downto 0);
constant uint1330_t_SLV_LEN : integer := 1330;
function uint1330_t_to_slv(x : uint1330_t) return std_logic_vector;
function slv_to_uint1330_t(x : std_logic_vector) return uint1330_t;
subtype int1330_t is signed(1329 downto 0);
constant int1330_t_SLV_LEN : integer := 1330;
function int1330_t_to_slv(x : int1330_t) return std_logic_vector;
function slv_to_int1330_t(x : std_logic_vector) return int1330_t;
subtype uint1331_t is unsigned(1330 downto 0);
constant uint1331_t_SLV_LEN : integer := 1331;
function uint1331_t_to_slv(x : uint1331_t) return std_logic_vector;
function slv_to_uint1331_t(x : std_logic_vector) return uint1331_t;
subtype int1331_t is signed(1330 downto 0);
constant int1331_t_SLV_LEN : integer := 1331;
function int1331_t_to_slv(x : int1331_t) return std_logic_vector;
function slv_to_int1331_t(x : std_logic_vector) return int1331_t;
subtype uint1332_t is unsigned(1331 downto 0);
constant uint1332_t_SLV_LEN : integer := 1332;
function uint1332_t_to_slv(x : uint1332_t) return std_logic_vector;
function slv_to_uint1332_t(x : std_logic_vector) return uint1332_t;
subtype int1332_t is signed(1331 downto 0);
constant int1332_t_SLV_LEN : integer := 1332;
function int1332_t_to_slv(x : int1332_t) return std_logic_vector;
function slv_to_int1332_t(x : std_logic_vector) return int1332_t;
subtype uint1333_t is unsigned(1332 downto 0);
constant uint1333_t_SLV_LEN : integer := 1333;
function uint1333_t_to_slv(x : uint1333_t) return std_logic_vector;
function slv_to_uint1333_t(x : std_logic_vector) return uint1333_t;
subtype int1333_t is signed(1332 downto 0);
constant int1333_t_SLV_LEN : integer := 1333;
function int1333_t_to_slv(x : int1333_t) return std_logic_vector;
function slv_to_int1333_t(x : std_logic_vector) return int1333_t;
subtype uint1334_t is unsigned(1333 downto 0);
constant uint1334_t_SLV_LEN : integer := 1334;
function uint1334_t_to_slv(x : uint1334_t) return std_logic_vector;
function slv_to_uint1334_t(x : std_logic_vector) return uint1334_t;
subtype int1334_t is signed(1333 downto 0);
constant int1334_t_SLV_LEN : integer := 1334;
function int1334_t_to_slv(x : int1334_t) return std_logic_vector;
function slv_to_int1334_t(x : std_logic_vector) return int1334_t;
subtype uint1335_t is unsigned(1334 downto 0);
constant uint1335_t_SLV_LEN : integer := 1335;
function uint1335_t_to_slv(x : uint1335_t) return std_logic_vector;
function slv_to_uint1335_t(x : std_logic_vector) return uint1335_t;
subtype int1335_t is signed(1334 downto 0);
constant int1335_t_SLV_LEN : integer := 1335;
function int1335_t_to_slv(x : int1335_t) return std_logic_vector;
function slv_to_int1335_t(x : std_logic_vector) return int1335_t;
subtype uint1336_t is unsigned(1335 downto 0);
constant uint1336_t_SLV_LEN : integer := 1336;
function uint1336_t_to_slv(x : uint1336_t) return std_logic_vector;
function slv_to_uint1336_t(x : std_logic_vector) return uint1336_t;
subtype int1336_t is signed(1335 downto 0);
constant int1336_t_SLV_LEN : integer := 1336;
function int1336_t_to_slv(x : int1336_t) return std_logic_vector;
function slv_to_int1336_t(x : std_logic_vector) return int1336_t;
subtype uint1337_t is unsigned(1336 downto 0);
constant uint1337_t_SLV_LEN : integer := 1337;
function uint1337_t_to_slv(x : uint1337_t) return std_logic_vector;
function slv_to_uint1337_t(x : std_logic_vector) return uint1337_t;
subtype int1337_t is signed(1336 downto 0);
constant int1337_t_SLV_LEN : integer := 1337;
function int1337_t_to_slv(x : int1337_t) return std_logic_vector;
function slv_to_int1337_t(x : std_logic_vector) return int1337_t;
subtype uint1338_t is unsigned(1337 downto 0);
constant uint1338_t_SLV_LEN : integer := 1338;
function uint1338_t_to_slv(x : uint1338_t) return std_logic_vector;
function slv_to_uint1338_t(x : std_logic_vector) return uint1338_t;
subtype int1338_t is signed(1337 downto 0);
constant int1338_t_SLV_LEN : integer := 1338;
function int1338_t_to_slv(x : int1338_t) return std_logic_vector;
function slv_to_int1338_t(x : std_logic_vector) return int1338_t;
subtype uint1339_t is unsigned(1338 downto 0);
constant uint1339_t_SLV_LEN : integer := 1339;
function uint1339_t_to_slv(x : uint1339_t) return std_logic_vector;
function slv_to_uint1339_t(x : std_logic_vector) return uint1339_t;
subtype int1339_t is signed(1338 downto 0);
constant int1339_t_SLV_LEN : integer := 1339;
function int1339_t_to_slv(x : int1339_t) return std_logic_vector;
function slv_to_int1339_t(x : std_logic_vector) return int1339_t;
subtype uint1340_t is unsigned(1339 downto 0);
constant uint1340_t_SLV_LEN : integer := 1340;
function uint1340_t_to_slv(x : uint1340_t) return std_logic_vector;
function slv_to_uint1340_t(x : std_logic_vector) return uint1340_t;
subtype int1340_t is signed(1339 downto 0);
constant int1340_t_SLV_LEN : integer := 1340;
function int1340_t_to_slv(x : int1340_t) return std_logic_vector;
function slv_to_int1340_t(x : std_logic_vector) return int1340_t;
subtype uint1341_t is unsigned(1340 downto 0);
constant uint1341_t_SLV_LEN : integer := 1341;
function uint1341_t_to_slv(x : uint1341_t) return std_logic_vector;
function slv_to_uint1341_t(x : std_logic_vector) return uint1341_t;
subtype int1341_t is signed(1340 downto 0);
constant int1341_t_SLV_LEN : integer := 1341;
function int1341_t_to_slv(x : int1341_t) return std_logic_vector;
function slv_to_int1341_t(x : std_logic_vector) return int1341_t;
subtype uint1342_t is unsigned(1341 downto 0);
constant uint1342_t_SLV_LEN : integer := 1342;
function uint1342_t_to_slv(x : uint1342_t) return std_logic_vector;
function slv_to_uint1342_t(x : std_logic_vector) return uint1342_t;
subtype int1342_t is signed(1341 downto 0);
constant int1342_t_SLV_LEN : integer := 1342;
function int1342_t_to_slv(x : int1342_t) return std_logic_vector;
function slv_to_int1342_t(x : std_logic_vector) return int1342_t;
subtype uint1343_t is unsigned(1342 downto 0);
constant uint1343_t_SLV_LEN : integer := 1343;
function uint1343_t_to_slv(x : uint1343_t) return std_logic_vector;
function slv_to_uint1343_t(x : std_logic_vector) return uint1343_t;
subtype int1343_t is signed(1342 downto 0);
constant int1343_t_SLV_LEN : integer := 1343;
function int1343_t_to_slv(x : int1343_t) return std_logic_vector;
function slv_to_int1343_t(x : std_logic_vector) return int1343_t;
subtype uint1344_t is unsigned(1343 downto 0);
constant uint1344_t_SLV_LEN : integer := 1344;
function uint1344_t_to_slv(x : uint1344_t) return std_logic_vector;
function slv_to_uint1344_t(x : std_logic_vector) return uint1344_t;
subtype int1344_t is signed(1343 downto 0);
constant int1344_t_SLV_LEN : integer := 1344;
function int1344_t_to_slv(x : int1344_t) return std_logic_vector;
function slv_to_int1344_t(x : std_logic_vector) return int1344_t;
subtype uint1345_t is unsigned(1344 downto 0);
constant uint1345_t_SLV_LEN : integer := 1345;
function uint1345_t_to_slv(x : uint1345_t) return std_logic_vector;
function slv_to_uint1345_t(x : std_logic_vector) return uint1345_t;
subtype int1345_t is signed(1344 downto 0);
constant int1345_t_SLV_LEN : integer := 1345;
function int1345_t_to_slv(x : int1345_t) return std_logic_vector;
function slv_to_int1345_t(x : std_logic_vector) return int1345_t;
subtype uint1346_t is unsigned(1345 downto 0);
constant uint1346_t_SLV_LEN : integer := 1346;
function uint1346_t_to_slv(x : uint1346_t) return std_logic_vector;
function slv_to_uint1346_t(x : std_logic_vector) return uint1346_t;
subtype int1346_t is signed(1345 downto 0);
constant int1346_t_SLV_LEN : integer := 1346;
function int1346_t_to_slv(x : int1346_t) return std_logic_vector;
function slv_to_int1346_t(x : std_logic_vector) return int1346_t;
subtype uint1347_t is unsigned(1346 downto 0);
constant uint1347_t_SLV_LEN : integer := 1347;
function uint1347_t_to_slv(x : uint1347_t) return std_logic_vector;
function slv_to_uint1347_t(x : std_logic_vector) return uint1347_t;
subtype int1347_t is signed(1346 downto 0);
constant int1347_t_SLV_LEN : integer := 1347;
function int1347_t_to_slv(x : int1347_t) return std_logic_vector;
function slv_to_int1347_t(x : std_logic_vector) return int1347_t;
subtype uint1348_t is unsigned(1347 downto 0);
constant uint1348_t_SLV_LEN : integer := 1348;
function uint1348_t_to_slv(x : uint1348_t) return std_logic_vector;
function slv_to_uint1348_t(x : std_logic_vector) return uint1348_t;
subtype int1348_t is signed(1347 downto 0);
constant int1348_t_SLV_LEN : integer := 1348;
function int1348_t_to_slv(x : int1348_t) return std_logic_vector;
function slv_to_int1348_t(x : std_logic_vector) return int1348_t;
subtype uint1349_t is unsigned(1348 downto 0);
constant uint1349_t_SLV_LEN : integer := 1349;
function uint1349_t_to_slv(x : uint1349_t) return std_logic_vector;
function slv_to_uint1349_t(x : std_logic_vector) return uint1349_t;
subtype int1349_t is signed(1348 downto 0);
constant int1349_t_SLV_LEN : integer := 1349;
function int1349_t_to_slv(x : int1349_t) return std_logic_vector;
function slv_to_int1349_t(x : std_logic_vector) return int1349_t;
subtype uint1350_t is unsigned(1349 downto 0);
constant uint1350_t_SLV_LEN : integer := 1350;
function uint1350_t_to_slv(x : uint1350_t) return std_logic_vector;
function slv_to_uint1350_t(x : std_logic_vector) return uint1350_t;
subtype int1350_t is signed(1349 downto 0);
constant int1350_t_SLV_LEN : integer := 1350;
function int1350_t_to_slv(x : int1350_t) return std_logic_vector;
function slv_to_int1350_t(x : std_logic_vector) return int1350_t;
subtype uint1351_t is unsigned(1350 downto 0);
constant uint1351_t_SLV_LEN : integer := 1351;
function uint1351_t_to_slv(x : uint1351_t) return std_logic_vector;
function slv_to_uint1351_t(x : std_logic_vector) return uint1351_t;
subtype int1351_t is signed(1350 downto 0);
constant int1351_t_SLV_LEN : integer := 1351;
function int1351_t_to_slv(x : int1351_t) return std_logic_vector;
function slv_to_int1351_t(x : std_logic_vector) return int1351_t;
subtype uint1352_t is unsigned(1351 downto 0);
constant uint1352_t_SLV_LEN : integer := 1352;
function uint1352_t_to_slv(x : uint1352_t) return std_logic_vector;
function slv_to_uint1352_t(x : std_logic_vector) return uint1352_t;
subtype int1352_t is signed(1351 downto 0);
constant int1352_t_SLV_LEN : integer := 1352;
function int1352_t_to_slv(x : int1352_t) return std_logic_vector;
function slv_to_int1352_t(x : std_logic_vector) return int1352_t;
subtype uint1353_t is unsigned(1352 downto 0);
constant uint1353_t_SLV_LEN : integer := 1353;
function uint1353_t_to_slv(x : uint1353_t) return std_logic_vector;
function slv_to_uint1353_t(x : std_logic_vector) return uint1353_t;
subtype int1353_t is signed(1352 downto 0);
constant int1353_t_SLV_LEN : integer := 1353;
function int1353_t_to_slv(x : int1353_t) return std_logic_vector;
function slv_to_int1353_t(x : std_logic_vector) return int1353_t;
subtype uint1354_t is unsigned(1353 downto 0);
constant uint1354_t_SLV_LEN : integer := 1354;
function uint1354_t_to_slv(x : uint1354_t) return std_logic_vector;
function slv_to_uint1354_t(x : std_logic_vector) return uint1354_t;
subtype int1354_t is signed(1353 downto 0);
constant int1354_t_SLV_LEN : integer := 1354;
function int1354_t_to_slv(x : int1354_t) return std_logic_vector;
function slv_to_int1354_t(x : std_logic_vector) return int1354_t;
subtype uint1355_t is unsigned(1354 downto 0);
constant uint1355_t_SLV_LEN : integer := 1355;
function uint1355_t_to_slv(x : uint1355_t) return std_logic_vector;
function slv_to_uint1355_t(x : std_logic_vector) return uint1355_t;
subtype int1355_t is signed(1354 downto 0);
constant int1355_t_SLV_LEN : integer := 1355;
function int1355_t_to_slv(x : int1355_t) return std_logic_vector;
function slv_to_int1355_t(x : std_logic_vector) return int1355_t;
subtype uint1356_t is unsigned(1355 downto 0);
constant uint1356_t_SLV_LEN : integer := 1356;
function uint1356_t_to_slv(x : uint1356_t) return std_logic_vector;
function slv_to_uint1356_t(x : std_logic_vector) return uint1356_t;
subtype int1356_t is signed(1355 downto 0);
constant int1356_t_SLV_LEN : integer := 1356;
function int1356_t_to_slv(x : int1356_t) return std_logic_vector;
function slv_to_int1356_t(x : std_logic_vector) return int1356_t;
subtype uint1357_t is unsigned(1356 downto 0);
constant uint1357_t_SLV_LEN : integer := 1357;
function uint1357_t_to_slv(x : uint1357_t) return std_logic_vector;
function slv_to_uint1357_t(x : std_logic_vector) return uint1357_t;
subtype int1357_t is signed(1356 downto 0);
constant int1357_t_SLV_LEN : integer := 1357;
function int1357_t_to_slv(x : int1357_t) return std_logic_vector;
function slv_to_int1357_t(x : std_logic_vector) return int1357_t;
subtype uint1358_t is unsigned(1357 downto 0);
constant uint1358_t_SLV_LEN : integer := 1358;
function uint1358_t_to_slv(x : uint1358_t) return std_logic_vector;
function slv_to_uint1358_t(x : std_logic_vector) return uint1358_t;
subtype int1358_t is signed(1357 downto 0);
constant int1358_t_SLV_LEN : integer := 1358;
function int1358_t_to_slv(x : int1358_t) return std_logic_vector;
function slv_to_int1358_t(x : std_logic_vector) return int1358_t;
subtype uint1359_t is unsigned(1358 downto 0);
constant uint1359_t_SLV_LEN : integer := 1359;
function uint1359_t_to_slv(x : uint1359_t) return std_logic_vector;
function slv_to_uint1359_t(x : std_logic_vector) return uint1359_t;
subtype int1359_t is signed(1358 downto 0);
constant int1359_t_SLV_LEN : integer := 1359;
function int1359_t_to_slv(x : int1359_t) return std_logic_vector;
function slv_to_int1359_t(x : std_logic_vector) return int1359_t;
subtype uint1360_t is unsigned(1359 downto 0);
constant uint1360_t_SLV_LEN : integer := 1360;
function uint1360_t_to_slv(x : uint1360_t) return std_logic_vector;
function slv_to_uint1360_t(x : std_logic_vector) return uint1360_t;
subtype int1360_t is signed(1359 downto 0);
constant int1360_t_SLV_LEN : integer := 1360;
function int1360_t_to_slv(x : int1360_t) return std_logic_vector;
function slv_to_int1360_t(x : std_logic_vector) return int1360_t;
subtype uint1361_t is unsigned(1360 downto 0);
constant uint1361_t_SLV_LEN : integer := 1361;
function uint1361_t_to_slv(x : uint1361_t) return std_logic_vector;
function slv_to_uint1361_t(x : std_logic_vector) return uint1361_t;
subtype int1361_t is signed(1360 downto 0);
constant int1361_t_SLV_LEN : integer := 1361;
function int1361_t_to_slv(x : int1361_t) return std_logic_vector;
function slv_to_int1361_t(x : std_logic_vector) return int1361_t;
subtype uint1362_t is unsigned(1361 downto 0);
constant uint1362_t_SLV_LEN : integer := 1362;
function uint1362_t_to_slv(x : uint1362_t) return std_logic_vector;
function slv_to_uint1362_t(x : std_logic_vector) return uint1362_t;
subtype int1362_t is signed(1361 downto 0);
constant int1362_t_SLV_LEN : integer := 1362;
function int1362_t_to_slv(x : int1362_t) return std_logic_vector;
function slv_to_int1362_t(x : std_logic_vector) return int1362_t;
subtype uint1363_t is unsigned(1362 downto 0);
constant uint1363_t_SLV_LEN : integer := 1363;
function uint1363_t_to_slv(x : uint1363_t) return std_logic_vector;
function slv_to_uint1363_t(x : std_logic_vector) return uint1363_t;
subtype int1363_t is signed(1362 downto 0);
constant int1363_t_SLV_LEN : integer := 1363;
function int1363_t_to_slv(x : int1363_t) return std_logic_vector;
function slv_to_int1363_t(x : std_logic_vector) return int1363_t;
subtype uint1364_t is unsigned(1363 downto 0);
constant uint1364_t_SLV_LEN : integer := 1364;
function uint1364_t_to_slv(x : uint1364_t) return std_logic_vector;
function slv_to_uint1364_t(x : std_logic_vector) return uint1364_t;
subtype int1364_t is signed(1363 downto 0);
constant int1364_t_SLV_LEN : integer := 1364;
function int1364_t_to_slv(x : int1364_t) return std_logic_vector;
function slv_to_int1364_t(x : std_logic_vector) return int1364_t;
subtype uint1365_t is unsigned(1364 downto 0);
constant uint1365_t_SLV_LEN : integer := 1365;
function uint1365_t_to_slv(x : uint1365_t) return std_logic_vector;
function slv_to_uint1365_t(x : std_logic_vector) return uint1365_t;
subtype int1365_t is signed(1364 downto 0);
constant int1365_t_SLV_LEN : integer := 1365;
function int1365_t_to_slv(x : int1365_t) return std_logic_vector;
function slv_to_int1365_t(x : std_logic_vector) return int1365_t;
subtype uint1366_t is unsigned(1365 downto 0);
constant uint1366_t_SLV_LEN : integer := 1366;
function uint1366_t_to_slv(x : uint1366_t) return std_logic_vector;
function slv_to_uint1366_t(x : std_logic_vector) return uint1366_t;
subtype int1366_t is signed(1365 downto 0);
constant int1366_t_SLV_LEN : integer := 1366;
function int1366_t_to_slv(x : int1366_t) return std_logic_vector;
function slv_to_int1366_t(x : std_logic_vector) return int1366_t;
subtype uint1367_t is unsigned(1366 downto 0);
constant uint1367_t_SLV_LEN : integer := 1367;
function uint1367_t_to_slv(x : uint1367_t) return std_logic_vector;
function slv_to_uint1367_t(x : std_logic_vector) return uint1367_t;
subtype int1367_t is signed(1366 downto 0);
constant int1367_t_SLV_LEN : integer := 1367;
function int1367_t_to_slv(x : int1367_t) return std_logic_vector;
function slv_to_int1367_t(x : std_logic_vector) return int1367_t;
subtype uint1368_t is unsigned(1367 downto 0);
constant uint1368_t_SLV_LEN : integer := 1368;
function uint1368_t_to_slv(x : uint1368_t) return std_logic_vector;
function slv_to_uint1368_t(x : std_logic_vector) return uint1368_t;
subtype int1368_t is signed(1367 downto 0);
constant int1368_t_SLV_LEN : integer := 1368;
function int1368_t_to_slv(x : int1368_t) return std_logic_vector;
function slv_to_int1368_t(x : std_logic_vector) return int1368_t;
subtype uint1369_t is unsigned(1368 downto 0);
constant uint1369_t_SLV_LEN : integer := 1369;
function uint1369_t_to_slv(x : uint1369_t) return std_logic_vector;
function slv_to_uint1369_t(x : std_logic_vector) return uint1369_t;
subtype int1369_t is signed(1368 downto 0);
constant int1369_t_SLV_LEN : integer := 1369;
function int1369_t_to_slv(x : int1369_t) return std_logic_vector;
function slv_to_int1369_t(x : std_logic_vector) return int1369_t;
subtype uint1370_t is unsigned(1369 downto 0);
constant uint1370_t_SLV_LEN : integer := 1370;
function uint1370_t_to_slv(x : uint1370_t) return std_logic_vector;
function slv_to_uint1370_t(x : std_logic_vector) return uint1370_t;
subtype int1370_t is signed(1369 downto 0);
constant int1370_t_SLV_LEN : integer := 1370;
function int1370_t_to_slv(x : int1370_t) return std_logic_vector;
function slv_to_int1370_t(x : std_logic_vector) return int1370_t;
subtype uint1371_t is unsigned(1370 downto 0);
constant uint1371_t_SLV_LEN : integer := 1371;
function uint1371_t_to_slv(x : uint1371_t) return std_logic_vector;
function slv_to_uint1371_t(x : std_logic_vector) return uint1371_t;
subtype int1371_t is signed(1370 downto 0);
constant int1371_t_SLV_LEN : integer := 1371;
function int1371_t_to_slv(x : int1371_t) return std_logic_vector;
function slv_to_int1371_t(x : std_logic_vector) return int1371_t;
subtype uint1372_t is unsigned(1371 downto 0);
constant uint1372_t_SLV_LEN : integer := 1372;
function uint1372_t_to_slv(x : uint1372_t) return std_logic_vector;
function slv_to_uint1372_t(x : std_logic_vector) return uint1372_t;
subtype int1372_t is signed(1371 downto 0);
constant int1372_t_SLV_LEN : integer := 1372;
function int1372_t_to_slv(x : int1372_t) return std_logic_vector;
function slv_to_int1372_t(x : std_logic_vector) return int1372_t;
subtype uint1373_t is unsigned(1372 downto 0);
constant uint1373_t_SLV_LEN : integer := 1373;
function uint1373_t_to_slv(x : uint1373_t) return std_logic_vector;
function slv_to_uint1373_t(x : std_logic_vector) return uint1373_t;
subtype int1373_t is signed(1372 downto 0);
constant int1373_t_SLV_LEN : integer := 1373;
function int1373_t_to_slv(x : int1373_t) return std_logic_vector;
function slv_to_int1373_t(x : std_logic_vector) return int1373_t;
subtype uint1374_t is unsigned(1373 downto 0);
constant uint1374_t_SLV_LEN : integer := 1374;
function uint1374_t_to_slv(x : uint1374_t) return std_logic_vector;
function slv_to_uint1374_t(x : std_logic_vector) return uint1374_t;
subtype int1374_t is signed(1373 downto 0);
constant int1374_t_SLV_LEN : integer := 1374;
function int1374_t_to_slv(x : int1374_t) return std_logic_vector;
function slv_to_int1374_t(x : std_logic_vector) return int1374_t;
subtype uint1375_t is unsigned(1374 downto 0);
constant uint1375_t_SLV_LEN : integer := 1375;
function uint1375_t_to_slv(x : uint1375_t) return std_logic_vector;
function slv_to_uint1375_t(x : std_logic_vector) return uint1375_t;
subtype int1375_t is signed(1374 downto 0);
constant int1375_t_SLV_LEN : integer := 1375;
function int1375_t_to_slv(x : int1375_t) return std_logic_vector;
function slv_to_int1375_t(x : std_logic_vector) return int1375_t;
subtype uint1376_t is unsigned(1375 downto 0);
constant uint1376_t_SLV_LEN : integer := 1376;
function uint1376_t_to_slv(x : uint1376_t) return std_logic_vector;
function slv_to_uint1376_t(x : std_logic_vector) return uint1376_t;
subtype int1376_t is signed(1375 downto 0);
constant int1376_t_SLV_LEN : integer := 1376;
function int1376_t_to_slv(x : int1376_t) return std_logic_vector;
function slv_to_int1376_t(x : std_logic_vector) return int1376_t;
subtype uint1377_t is unsigned(1376 downto 0);
constant uint1377_t_SLV_LEN : integer := 1377;
function uint1377_t_to_slv(x : uint1377_t) return std_logic_vector;
function slv_to_uint1377_t(x : std_logic_vector) return uint1377_t;
subtype int1377_t is signed(1376 downto 0);
constant int1377_t_SLV_LEN : integer := 1377;
function int1377_t_to_slv(x : int1377_t) return std_logic_vector;
function slv_to_int1377_t(x : std_logic_vector) return int1377_t;
subtype uint1378_t is unsigned(1377 downto 0);
constant uint1378_t_SLV_LEN : integer := 1378;
function uint1378_t_to_slv(x : uint1378_t) return std_logic_vector;
function slv_to_uint1378_t(x : std_logic_vector) return uint1378_t;
subtype int1378_t is signed(1377 downto 0);
constant int1378_t_SLV_LEN : integer := 1378;
function int1378_t_to_slv(x : int1378_t) return std_logic_vector;
function slv_to_int1378_t(x : std_logic_vector) return int1378_t;
subtype uint1379_t is unsigned(1378 downto 0);
constant uint1379_t_SLV_LEN : integer := 1379;
function uint1379_t_to_slv(x : uint1379_t) return std_logic_vector;
function slv_to_uint1379_t(x : std_logic_vector) return uint1379_t;
subtype int1379_t is signed(1378 downto 0);
constant int1379_t_SLV_LEN : integer := 1379;
function int1379_t_to_slv(x : int1379_t) return std_logic_vector;
function slv_to_int1379_t(x : std_logic_vector) return int1379_t;
subtype uint1380_t is unsigned(1379 downto 0);
constant uint1380_t_SLV_LEN : integer := 1380;
function uint1380_t_to_slv(x : uint1380_t) return std_logic_vector;
function slv_to_uint1380_t(x : std_logic_vector) return uint1380_t;
subtype int1380_t is signed(1379 downto 0);
constant int1380_t_SLV_LEN : integer := 1380;
function int1380_t_to_slv(x : int1380_t) return std_logic_vector;
function slv_to_int1380_t(x : std_logic_vector) return int1380_t;
subtype uint1381_t is unsigned(1380 downto 0);
constant uint1381_t_SLV_LEN : integer := 1381;
function uint1381_t_to_slv(x : uint1381_t) return std_logic_vector;
function slv_to_uint1381_t(x : std_logic_vector) return uint1381_t;
subtype int1381_t is signed(1380 downto 0);
constant int1381_t_SLV_LEN : integer := 1381;
function int1381_t_to_slv(x : int1381_t) return std_logic_vector;
function slv_to_int1381_t(x : std_logic_vector) return int1381_t;
subtype uint1382_t is unsigned(1381 downto 0);
constant uint1382_t_SLV_LEN : integer := 1382;
function uint1382_t_to_slv(x : uint1382_t) return std_logic_vector;
function slv_to_uint1382_t(x : std_logic_vector) return uint1382_t;
subtype int1382_t is signed(1381 downto 0);
constant int1382_t_SLV_LEN : integer := 1382;
function int1382_t_to_slv(x : int1382_t) return std_logic_vector;
function slv_to_int1382_t(x : std_logic_vector) return int1382_t;
subtype uint1383_t is unsigned(1382 downto 0);
constant uint1383_t_SLV_LEN : integer := 1383;
function uint1383_t_to_slv(x : uint1383_t) return std_logic_vector;
function slv_to_uint1383_t(x : std_logic_vector) return uint1383_t;
subtype int1383_t is signed(1382 downto 0);
constant int1383_t_SLV_LEN : integer := 1383;
function int1383_t_to_slv(x : int1383_t) return std_logic_vector;
function slv_to_int1383_t(x : std_logic_vector) return int1383_t;
subtype uint1384_t is unsigned(1383 downto 0);
constant uint1384_t_SLV_LEN : integer := 1384;
function uint1384_t_to_slv(x : uint1384_t) return std_logic_vector;
function slv_to_uint1384_t(x : std_logic_vector) return uint1384_t;
subtype int1384_t is signed(1383 downto 0);
constant int1384_t_SLV_LEN : integer := 1384;
function int1384_t_to_slv(x : int1384_t) return std_logic_vector;
function slv_to_int1384_t(x : std_logic_vector) return int1384_t;
subtype uint1385_t is unsigned(1384 downto 0);
constant uint1385_t_SLV_LEN : integer := 1385;
function uint1385_t_to_slv(x : uint1385_t) return std_logic_vector;
function slv_to_uint1385_t(x : std_logic_vector) return uint1385_t;
subtype int1385_t is signed(1384 downto 0);
constant int1385_t_SLV_LEN : integer := 1385;
function int1385_t_to_slv(x : int1385_t) return std_logic_vector;
function slv_to_int1385_t(x : std_logic_vector) return int1385_t;
subtype uint1386_t is unsigned(1385 downto 0);
constant uint1386_t_SLV_LEN : integer := 1386;
function uint1386_t_to_slv(x : uint1386_t) return std_logic_vector;
function slv_to_uint1386_t(x : std_logic_vector) return uint1386_t;
subtype int1386_t is signed(1385 downto 0);
constant int1386_t_SLV_LEN : integer := 1386;
function int1386_t_to_slv(x : int1386_t) return std_logic_vector;
function slv_to_int1386_t(x : std_logic_vector) return int1386_t;
subtype uint1387_t is unsigned(1386 downto 0);
constant uint1387_t_SLV_LEN : integer := 1387;
function uint1387_t_to_slv(x : uint1387_t) return std_logic_vector;
function slv_to_uint1387_t(x : std_logic_vector) return uint1387_t;
subtype int1387_t is signed(1386 downto 0);
constant int1387_t_SLV_LEN : integer := 1387;
function int1387_t_to_slv(x : int1387_t) return std_logic_vector;
function slv_to_int1387_t(x : std_logic_vector) return int1387_t;
subtype uint1388_t is unsigned(1387 downto 0);
constant uint1388_t_SLV_LEN : integer := 1388;
function uint1388_t_to_slv(x : uint1388_t) return std_logic_vector;
function slv_to_uint1388_t(x : std_logic_vector) return uint1388_t;
subtype int1388_t is signed(1387 downto 0);
constant int1388_t_SLV_LEN : integer := 1388;
function int1388_t_to_slv(x : int1388_t) return std_logic_vector;
function slv_to_int1388_t(x : std_logic_vector) return int1388_t;
subtype uint1389_t is unsigned(1388 downto 0);
constant uint1389_t_SLV_LEN : integer := 1389;
function uint1389_t_to_slv(x : uint1389_t) return std_logic_vector;
function slv_to_uint1389_t(x : std_logic_vector) return uint1389_t;
subtype int1389_t is signed(1388 downto 0);
constant int1389_t_SLV_LEN : integer := 1389;
function int1389_t_to_slv(x : int1389_t) return std_logic_vector;
function slv_to_int1389_t(x : std_logic_vector) return int1389_t;
subtype uint1390_t is unsigned(1389 downto 0);
constant uint1390_t_SLV_LEN : integer := 1390;
function uint1390_t_to_slv(x : uint1390_t) return std_logic_vector;
function slv_to_uint1390_t(x : std_logic_vector) return uint1390_t;
subtype int1390_t is signed(1389 downto 0);
constant int1390_t_SLV_LEN : integer := 1390;
function int1390_t_to_slv(x : int1390_t) return std_logic_vector;
function slv_to_int1390_t(x : std_logic_vector) return int1390_t;
subtype uint1391_t is unsigned(1390 downto 0);
constant uint1391_t_SLV_LEN : integer := 1391;
function uint1391_t_to_slv(x : uint1391_t) return std_logic_vector;
function slv_to_uint1391_t(x : std_logic_vector) return uint1391_t;
subtype int1391_t is signed(1390 downto 0);
constant int1391_t_SLV_LEN : integer := 1391;
function int1391_t_to_slv(x : int1391_t) return std_logic_vector;
function slv_to_int1391_t(x : std_logic_vector) return int1391_t;
subtype uint1392_t is unsigned(1391 downto 0);
constant uint1392_t_SLV_LEN : integer := 1392;
function uint1392_t_to_slv(x : uint1392_t) return std_logic_vector;
function slv_to_uint1392_t(x : std_logic_vector) return uint1392_t;
subtype int1392_t is signed(1391 downto 0);
constant int1392_t_SLV_LEN : integer := 1392;
function int1392_t_to_slv(x : int1392_t) return std_logic_vector;
function slv_to_int1392_t(x : std_logic_vector) return int1392_t;
subtype uint1393_t is unsigned(1392 downto 0);
constant uint1393_t_SLV_LEN : integer := 1393;
function uint1393_t_to_slv(x : uint1393_t) return std_logic_vector;
function slv_to_uint1393_t(x : std_logic_vector) return uint1393_t;
subtype int1393_t is signed(1392 downto 0);
constant int1393_t_SLV_LEN : integer := 1393;
function int1393_t_to_slv(x : int1393_t) return std_logic_vector;
function slv_to_int1393_t(x : std_logic_vector) return int1393_t;
subtype uint1394_t is unsigned(1393 downto 0);
constant uint1394_t_SLV_LEN : integer := 1394;
function uint1394_t_to_slv(x : uint1394_t) return std_logic_vector;
function slv_to_uint1394_t(x : std_logic_vector) return uint1394_t;
subtype int1394_t is signed(1393 downto 0);
constant int1394_t_SLV_LEN : integer := 1394;
function int1394_t_to_slv(x : int1394_t) return std_logic_vector;
function slv_to_int1394_t(x : std_logic_vector) return int1394_t;
subtype uint1395_t is unsigned(1394 downto 0);
constant uint1395_t_SLV_LEN : integer := 1395;
function uint1395_t_to_slv(x : uint1395_t) return std_logic_vector;
function slv_to_uint1395_t(x : std_logic_vector) return uint1395_t;
subtype int1395_t is signed(1394 downto 0);
constant int1395_t_SLV_LEN : integer := 1395;
function int1395_t_to_slv(x : int1395_t) return std_logic_vector;
function slv_to_int1395_t(x : std_logic_vector) return int1395_t;
subtype uint1396_t is unsigned(1395 downto 0);
constant uint1396_t_SLV_LEN : integer := 1396;
function uint1396_t_to_slv(x : uint1396_t) return std_logic_vector;
function slv_to_uint1396_t(x : std_logic_vector) return uint1396_t;
subtype int1396_t is signed(1395 downto 0);
constant int1396_t_SLV_LEN : integer := 1396;
function int1396_t_to_slv(x : int1396_t) return std_logic_vector;
function slv_to_int1396_t(x : std_logic_vector) return int1396_t;
subtype uint1397_t is unsigned(1396 downto 0);
constant uint1397_t_SLV_LEN : integer := 1397;
function uint1397_t_to_slv(x : uint1397_t) return std_logic_vector;
function slv_to_uint1397_t(x : std_logic_vector) return uint1397_t;
subtype int1397_t is signed(1396 downto 0);
constant int1397_t_SLV_LEN : integer := 1397;
function int1397_t_to_slv(x : int1397_t) return std_logic_vector;
function slv_to_int1397_t(x : std_logic_vector) return int1397_t;
subtype uint1398_t is unsigned(1397 downto 0);
constant uint1398_t_SLV_LEN : integer := 1398;
function uint1398_t_to_slv(x : uint1398_t) return std_logic_vector;
function slv_to_uint1398_t(x : std_logic_vector) return uint1398_t;
subtype int1398_t is signed(1397 downto 0);
constant int1398_t_SLV_LEN : integer := 1398;
function int1398_t_to_slv(x : int1398_t) return std_logic_vector;
function slv_to_int1398_t(x : std_logic_vector) return int1398_t;
subtype uint1399_t is unsigned(1398 downto 0);
constant uint1399_t_SLV_LEN : integer := 1399;
function uint1399_t_to_slv(x : uint1399_t) return std_logic_vector;
function slv_to_uint1399_t(x : std_logic_vector) return uint1399_t;
subtype int1399_t is signed(1398 downto 0);
constant int1399_t_SLV_LEN : integer := 1399;
function int1399_t_to_slv(x : int1399_t) return std_logic_vector;
function slv_to_int1399_t(x : std_logic_vector) return int1399_t;
subtype uint1400_t is unsigned(1399 downto 0);
constant uint1400_t_SLV_LEN : integer := 1400;
function uint1400_t_to_slv(x : uint1400_t) return std_logic_vector;
function slv_to_uint1400_t(x : std_logic_vector) return uint1400_t;
subtype int1400_t is signed(1399 downto 0);
constant int1400_t_SLV_LEN : integer := 1400;
function int1400_t_to_slv(x : int1400_t) return std_logic_vector;
function slv_to_int1400_t(x : std_logic_vector) return int1400_t;
subtype uint1401_t is unsigned(1400 downto 0);
constant uint1401_t_SLV_LEN : integer := 1401;
function uint1401_t_to_slv(x : uint1401_t) return std_logic_vector;
function slv_to_uint1401_t(x : std_logic_vector) return uint1401_t;
subtype int1401_t is signed(1400 downto 0);
constant int1401_t_SLV_LEN : integer := 1401;
function int1401_t_to_slv(x : int1401_t) return std_logic_vector;
function slv_to_int1401_t(x : std_logic_vector) return int1401_t;
subtype uint1402_t is unsigned(1401 downto 0);
constant uint1402_t_SLV_LEN : integer := 1402;
function uint1402_t_to_slv(x : uint1402_t) return std_logic_vector;
function slv_to_uint1402_t(x : std_logic_vector) return uint1402_t;
subtype int1402_t is signed(1401 downto 0);
constant int1402_t_SLV_LEN : integer := 1402;
function int1402_t_to_slv(x : int1402_t) return std_logic_vector;
function slv_to_int1402_t(x : std_logic_vector) return int1402_t;
subtype uint1403_t is unsigned(1402 downto 0);
constant uint1403_t_SLV_LEN : integer := 1403;
function uint1403_t_to_slv(x : uint1403_t) return std_logic_vector;
function slv_to_uint1403_t(x : std_logic_vector) return uint1403_t;
subtype int1403_t is signed(1402 downto 0);
constant int1403_t_SLV_LEN : integer := 1403;
function int1403_t_to_slv(x : int1403_t) return std_logic_vector;
function slv_to_int1403_t(x : std_logic_vector) return int1403_t;
subtype uint1404_t is unsigned(1403 downto 0);
constant uint1404_t_SLV_LEN : integer := 1404;
function uint1404_t_to_slv(x : uint1404_t) return std_logic_vector;
function slv_to_uint1404_t(x : std_logic_vector) return uint1404_t;
subtype int1404_t is signed(1403 downto 0);
constant int1404_t_SLV_LEN : integer := 1404;
function int1404_t_to_slv(x : int1404_t) return std_logic_vector;
function slv_to_int1404_t(x : std_logic_vector) return int1404_t;
subtype uint1405_t is unsigned(1404 downto 0);
constant uint1405_t_SLV_LEN : integer := 1405;
function uint1405_t_to_slv(x : uint1405_t) return std_logic_vector;
function slv_to_uint1405_t(x : std_logic_vector) return uint1405_t;
subtype int1405_t is signed(1404 downto 0);
constant int1405_t_SLV_LEN : integer := 1405;
function int1405_t_to_slv(x : int1405_t) return std_logic_vector;
function slv_to_int1405_t(x : std_logic_vector) return int1405_t;
subtype uint1406_t is unsigned(1405 downto 0);
constant uint1406_t_SLV_LEN : integer := 1406;
function uint1406_t_to_slv(x : uint1406_t) return std_logic_vector;
function slv_to_uint1406_t(x : std_logic_vector) return uint1406_t;
subtype int1406_t is signed(1405 downto 0);
constant int1406_t_SLV_LEN : integer := 1406;
function int1406_t_to_slv(x : int1406_t) return std_logic_vector;
function slv_to_int1406_t(x : std_logic_vector) return int1406_t;
subtype uint1407_t is unsigned(1406 downto 0);
constant uint1407_t_SLV_LEN : integer := 1407;
function uint1407_t_to_slv(x : uint1407_t) return std_logic_vector;
function slv_to_uint1407_t(x : std_logic_vector) return uint1407_t;
subtype int1407_t is signed(1406 downto 0);
constant int1407_t_SLV_LEN : integer := 1407;
function int1407_t_to_slv(x : int1407_t) return std_logic_vector;
function slv_to_int1407_t(x : std_logic_vector) return int1407_t;
subtype uint1408_t is unsigned(1407 downto 0);
constant uint1408_t_SLV_LEN : integer := 1408;
function uint1408_t_to_slv(x : uint1408_t) return std_logic_vector;
function slv_to_uint1408_t(x : std_logic_vector) return uint1408_t;
subtype int1408_t is signed(1407 downto 0);
constant int1408_t_SLV_LEN : integer := 1408;
function int1408_t_to_slv(x : int1408_t) return std_logic_vector;
function slv_to_int1408_t(x : std_logic_vector) return int1408_t;
subtype uint1409_t is unsigned(1408 downto 0);
constant uint1409_t_SLV_LEN : integer := 1409;
function uint1409_t_to_slv(x : uint1409_t) return std_logic_vector;
function slv_to_uint1409_t(x : std_logic_vector) return uint1409_t;
subtype int1409_t is signed(1408 downto 0);
constant int1409_t_SLV_LEN : integer := 1409;
function int1409_t_to_slv(x : int1409_t) return std_logic_vector;
function slv_to_int1409_t(x : std_logic_vector) return int1409_t;
subtype uint1410_t is unsigned(1409 downto 0);
constant uint1410_t_SLV_LEN : integer := 1410;
function uint1410_t_to_slv(x : uint1410_t) return std_logic_vector;
function slv_to_uint1410_t(x : std_logic_vector) return uint1410_t;
subtype int1410_t is signed(1409 downto 0);
constant int1410_t_SLV_LEN : integer := 1410;
function int1410_t_to_slv(x : int1410_t) return std_logic_vector;
function slv_to_int1410_t(x : std_logic_vector) return int1410_t;
subtype uint1411_t is unsigned(1410 downto 0);
constant uint1411_t_SLV_LEN : integer := 1411;
function uint1411_t_to_slv(x : uint1411_t) return std_logic_vector;
function slv_to_uint1411_t(x : std_logic_vector) return uint1411_t;
subtype int1411_t is signed(1410 downto 0);
constant int1411_t_SLV_LEN : integer := 1411;
function int1411_t_to_slv(x : int1411_t) return std_logic_vector;
function slv_to_int1411_t(x : std_logic_vector) return int1411_t;
subtype uint1412_t is unsigned(1411 downto 0);
constant uint1412_t_SLV_LEN : integer := 1412;
function uint1412_t_to_slv(x : uint1412_t) return std_logic_vector;
function slv_to_uint1412_t(x : std_logic_vector) return uint1412_t;
subtype int1412_t is signed(1411 downto 0);
constant int1412_t_SLV_LEN : integer := 1412;
function int1412_t_to_slv(x : int1412_t) return std_logic_vector;
function slv_to_int1412_t(x : std_logic_vector) return int1412_t;
subtype uint1413_t is unsigned(1412 downto 0);
constant uint1413_t_SLV_LEN : integer := 1413;
function uint1413_t_to_slv(x : uint1413_t) return std_logic_vector;
function slv_to_uint1413_t(x : std_logic_vector) return uint1413_t;
subtype int1413_t is signed(1412 downto 0);
constant int1413_t_SLV_LEN : integer := 1413;
function int1413_t_to_slv(x : int1413_t) return std_logic_vector;
function slv_to_int1413_t(x : std_logic_vector) return int1413_t;
subtype uint1414_t is unsigned(1413 downto 0);
constant uint1414_t_SLV_LEN : integer := 1414;
function uint1414_t_to_slv(x : uint1414_t) return std_logic_vector;
function slv_to_uint1414_t(x : std_logic_vector) return uint1414_t;
subtype int1414_t is signed(1413 downto 0);
constant int1414_t_SLV_LEN : integer := 1414;
function int1414_t_to_slv(x : int1414_t) return std_logic_vector;
function slv_to_int1414_t(x : std_logic_vector) return int1414_t;
subtype uint1415_t is unsigned(1414 downto 0);
constant uint1415_t_SLV_LEN : integer := 1415;
function uint1415_t_to_slv(x : uint1415_t) return std_logic_vector;
function slv_to_uint1415_t(x : std_logic_vector) return uint1415_t;
subtype int1415_t is signed(1414 downto 0);
constant int1415_t_SLV_LEN : integer := 1415;
function int1415_t_to_slv(x : int1415_t) return std_logic_vector;
function slv_to_int1415_t(x : std_logic_vector) return int1415_t;
subtype uint1416_t is unsigned(1415 downto 0);
constant uint1416_t_SLV_LEN : integer := 1416;
function uint1416_t_to_slv(x : uint1416_t) return std_logic_vector;
function slv_to_uint1416_t(x : std_logic_vector) return uint1416_t;
subtype int1416_t is signed(1415 downto 0);
constant int1416_t_SLV_LEN : integer := 1416;
function int1416_t_to_slv(x : int1416_t) return std_logic_vector;
function slv_to_int1416_t(x : std_logic_vector) return int1416_t;
subtype uint1417_t is unsigned(1416 downto 0);
constant uint1417_t_SLV_LEN : integer := 1417;
function uint1417_t_to_slv(x : uint1417_t) return std_logic_vector;
function slv_to_uint1417_t(x : std_logic_vector) return uint1417_t;
subtype int1417_t is signed(1416 downto 0);
constant int1417_t_SLV_LEN : integer := 1417;
function int1417_t_to_slv(x : int1417_t) return std_logic_vector;
function slv_to_int1417_t(x : std_logic_vector) return int1417_t;
subtype uint1418_t is unsigned(1417 downto 0);
constant uint1418_t_SLV_LEN : integer := 1418;
function uint1418_t_to_slv(x : uint1418_t) return std_logic_vector;
function slv_to_uint1418_t(x : std_logic_vector) return uint1418_t;
subtype int1418_t is signed(1417 downto 0);
constant int1418_t_SLV_LEN : integer := 1418;
function int1418_t_to_slv(x : int1418_t) return std_logic_vector;
function slv_to_int1418_t(x : std_logic_vector) return int1418_t;
subtype uint1419_t is unsigned(1418 downto 0);
constant uint1419_t_SLV_LEN : integer := 1419;
function uint1419_t_to_slv(x : uint1419_t) return std_logic_vector;
function slv_to_uint1419_t(x : std_logic_vector) return uint1419_t;
subtype int1419_t is signed(1418 downto 0);
constant int1419_t_SLV_LEN : integer := 1419;
function int1419_t_to_slv(x : int1419_t) return std_logic_vector;
function slv_to_int1419_t(x : std_logic_vector) return int1419_t;
subtype uint1420_t is unsigned(1419 downto 0);
constant uint1420_t_SLV_LEN : integer := 1420;
function uint1420_t_to_slv(x : uint1420_t) return std_logic_vector;
function slv_to_uint1420_t(x : std_logic_vector) return uint1420_t;
subtype int1420_t is signed(1419 downto 0);
constant int1420_t_SLV_LEN : integer := 1420;
function int1420_t_to_slv(x : int1420_t) return std_logic_vector;
function slv_to_int1420_t(x : std_logic_vector) return int1420_t;
subtype uint1421_t is unsigned(1420 downto 0);
constant uint1421_t_SLV_LEN : integer := 1421;
function uint1421_t_to_slv(x : uint1421_t) return std_logic_vector;
function slv_to_uint1421_t(x : std_logic_vector) return uint1421_t;
subtype int1421_t is signed(1420 downto 0);
constant int1421_t_SLV_LEN : integer := 1421;
function int1421_t_to_slv(x : int1421_t) return std_logic_vector;
function slv_to_int1421_t(x : std_logic_vector) return int1421_t;
subtype uint1422_t is unsigned(1421 downto 0);
constant uint1422_t_SLV_LEN : integer := 1422;
function uint1422_t_to_slv(x : uint1422_t) return std_logic_vector;
function slv_to_uint1422_t(x : std_logic_vector) return uint1422_t;
subtype int1422_t is signed(1421 downto 0);
constant int1422_t_SLV_LEN : integer := 1422;
function int1422_t_to_slv(x : int1422_t) return std_logic_vector;
function slv_to_int1422_t(x : std_logic_vector) return int1422_t;
subtype uint1423_t is unsigned(1422 downto 0);
constant uint1423_t_SLV_LEN : integer := 1423;
function uint1423_t_to_slv(x : uint1423_t) return std_logic_vector;
function slv_to_uint1423_t(x : std_logic_vector) return uint1423_t;
subtype int1423_t is signed(1422 downto 0);
constant int1423_t_SLV_LEN : integer := 1423;
function int1423_t_to_slv(x : int1423_t) return std_logic_vector;
function slv_to_int1423_t(x : std_logic_vector) return int1423_t;
subtype uint1424_t is unsigned(1423 downto 0);
constant uint1424_t_SLV_LEN : integer := 1424;
function uint1424_t_to_slv(x : uint1424_t) return std_logic_vector;
function slv_to_uint1424_t(x : std_logic_vector) return uint1424_t;
subtype int1424_t is signed(1423 downto 0);
constant int1424_t_SLV_LEN : integer := 1424;
function int1424_t_to_slv(x : int1424_t) return std_logic_vector;
function slv_to_int1424_t(x : std_logic_vector) return int1424_t;
subtype uint1425_t is unsigned(1424 downto 0);
constant uint1425_t_SLV_LEN : integer := 1425;
function uint1425_t_to_slv(x : uint1425_t) return std_logic_vector;
function slv_to_uint1425_t(x : std_logic_vector) return uint1425_t;
subtype int1425_t is signed(1424 downto 0);
constant int1425_t_SLV_LEN : integer := 1425;
function int1425_t_to_slv(x : int1425_t) return std_logic_vector;
function slv_to_int1425_t(x : std_logic_vector) return int1425_t;
subtype uint1426_t is unsigned(1425 downto 0);
constant uint1426_t_SLV_LEN : integer := 1426;
function uint1426_t_to_slv(x : uint1426_t) return std_logic_vector;
function slv_to_uint1426_t(x : std_logic_vector) return uint1426_t;
subtype int1426_t is signed(1425 downto 0);
constant int1426_t_SLV_LEN : integer := 1426;
function int1426_t_to_slv(x : int1426_t) return std_logic_vector;
function slv_to_int1426_t(x : std_logic_vector) return int1426_t;
subtype uint1427_t is unsigned(1426 downto 0);
constant uint1427_t_SLV_LEN : integer := 1427;
function uint1427_t_to_slv(x : uint1427_t) return std_logic_vector;
function slv_to_uint1427_t(x : std_logic_vector) return uint1427_t;
subtype int1427_t is signed(1426 downto 0);
constant int1427_t_SLV_LEN : integer := 1427;
function int1427_t_to_slv(x : int1427_t) return std_logic_vector;
function slv_to_int1427_t(x : std_logic_vector) return int1427_t;
subtype uint1428_t is unsigned(1427 downto 0);
constant uint1428_t_SLV_LEN : integer := 1428;
function uint1428_t_to_slv(x : uint1428_t) return std_logic_vector;
function slv_to_uint1428_t(x : std_logic_vector) return uint1428_t;
subtype int1428_t is signed(1427 downto 0);
constant int1428_t_SLV_LEN : integer := 1428;
function int1428_t_to_slv(x : int1428_t) return std_logic_vector;
function slv_to_int1428_t(x : std_logic_vector) return int1428_t;
subtype uint1429_t is unsigned(1428 downto 0);
constant uint1429_t_SLV_LEN : integer := 1429;
function uint1429_t_to_slv(x : uint1429_t) return std_logic_vector;
function slv_to_uint1429_t(x : std_logic_vector) return uint1429_t;
subtype int1429_t is signed(1428 downto 0);
constant int1429_t_SLV_LEN : integer := 1429;
function int1429_t_to_slv(x : int1429_t) return std_logic_vector;
function slv_to_int1429_t(x : std_logic_vector) return int1429_t;
subtype uint1430_t is unsigned(1429 downto 0);
constant uint1430_t_SLV_LEN : integer := 1430;
function uint1430_t_to_slv(x : uint1430_t) return std_logic_vector;
function slv_to_uint1430_t(x : std_logic_vector) return uint1430_t;
subtype int1430_t is signed(1429 downto 0);
constant int1430_t_SLV_LEN : integer := 1430;
function int1430_t_to_slv(x : int1430_t) return std_logic_vector;
function slv_to_int1430_t(x : std_logic_vector) return int1430_t;
subtype uint1431_t is unsigned(1430 downto 0);
constant uint1431_t_SLV_LEN : integer := 1431;
function uint1431_t_to_slv(x : uint1431_t) return std_logic_vector;
function slv_to_uint1431_t(x : std_logic_vector) return uint1431_t;
subtype int1431_t is signed(1430 downto 0);
constant int1431_t_SLV_LEN : integer := 1431;
function int1431_t_to_slv(x : int1431_t) return std_logic_vector;
function slv_to_int1431_t(x : std_logic_vector) return int1431_t;
subtype uint1432_t is unsigned(1431 downto 0);
constant uint1432_t_SLV_LEN : integer := 1432;
function uint1432_t_to_slv(x : uint1432_t) return std_logic_vector;
function slv_to_uint1432_t(x : std_logic_vector) return uint1432_t;
subtype int1432_t is signed(1431 downto 0);
constant int1432_t_SLV_LEN : integer := 1432;
function int1432_t_to_slv(x : int1432_t) return std_logic_vector;
function slv_to_int1432_t(x : std_logic_vector) return int1432_t;
subtype uint1433_t is unsigned(1432 downto 0);
constant uint1433_t_SLV_LEN : integer := 1433;
function uint1433_t_to_slv(x : uint1433_t) return std_logic_vector;
function slv_to_uint1433_t(x : std_logic_vector) return uint1433_t;
subtype int1433_t is signed(1432 downto 0);
constant int1433_t_SLV_LEN : integer := 1433;
function int1433_t_to_slv(x : int1433_t) return std_logic_vector;
function slv_to_int1433_t(x : std_logic_vector) return int1433_t;
subtype uint1434_t is unsigned(1433 downto 0);
constant uint1434_t_SLV_LEN : integer := 1434;
function uint1434_t_to_slv(x : uint1434_t) return std_logic_vector;
function slv_to_uint1434_t(x : std_logic_vector) return uint1434_t;
subtype int1434_t is signed(1433 downto 0);
constant int1434_t_SLV_LEN : integer := 1434;
function int1434_t_to_slv(x : int1434_t) return std_logic_vector;
function slv_to_int1434_t(x : std_logic_vector) return int1434_t;
subtype uint1435_t is unsigned(1434 downto 0);
constant uint1435_t_SLV_LEN : integer := 1435;
function uint1435_t_to_slv(x : uint1435_t) return std_logic_vector;
function slv_to_uint1435_t(x : std_logic_vector) return uint1435_t;
subtype int1435_t is signed(1434 downto 0);
constant int1435_t_SLV_LEN : integer := 1435;
function int1435_t_to_slv(x : int1435_t) return std_logic_vector;
function slv_to_int1435_t(x : std_logic_vector) return int1435_t;
subtype uint1436_t is unsigned(1435 downto 0);
constant uint1436_t_SLV_LEN : integer := 1436;
function uint1436_t_to_slv(x : uint1436_t) return std_logic_vector;
function slv_to_uint1436_t(x : std_logic_vector) return uint1436_t;
subtype int1436_t is signed(1435 downto 0);
constant int1436_t_SLV_LEN : integer := 1436;
function int1436_t_to_slv(x : int1436_t) return std_logic_vector;
function slv_to_int1436_t(x : std_logic_vector) return int1436_t;
subtype uint1437_t is unsigned(1436 downto 0);
constant uint1437_t_SLV_LEN : integer := 1437;
function uint1437_t_to_slv(x : uint1437_t) return std_logic_vector;
function slv_to_uint1437_t(x : std_logic_vector) return uint1437_t;
subtype int1437_t is signed(1436 downto 0);
constant int1437_t_SLV_LEN : integer := 1437;
function int1437_t_to_slv(x : int1437_t) return std_logic_vector;
function slv_to_int1437_t(x : std_logic_vector) return int1437_t;
subtype uint1438_t is unsigned(1437 downto 0);
constant uint1438_t_SLV_LEN : integer := 1438;
function uint1438_t_to_slv(x : uint1438_t) return std_logic_vector;
function slv_to_uint1438_t(x : std_logic_vector) return uint1438_t;
subtype int1438_t is signed(1437 downto 0);
constant int1438_t_SLV_LEN : integer := 1438;
function int1438_t_to_slv(x : int1438_t) return std_logic_vector;
function slv_to_int1438_t(x : std_logic_vector) return int1438_t;
subtype uint1439_t is unsigned(1438 downto 0);
constant uint1439_t_SLV_LEN : integer := 1439;
function uint1439_t_to_slv(x : uint1439_t) return std_logic_vector;
function slv_to_uint1439_t(x : std_logic_vector) return uint1439_t;
subtype int1439_t is signed(1438 downto 0);
constant int1439_t_SLV_LEN : integer := 1439;
function int1439_t_to_slv(x : int1439_t) return std_logic_vector;
function slv_to_int1439_t(x : std_logic_vector) return int1439_t;
subtype uint1440_t is unsigned(1439 downto 0);
constant uint1440_t_SLV_LEN : integer := 1440;
function uint1440_t_to_slv(x : uint1440_t) return std_logic_vector;
function slv_to_uint1440_t(x : std_logic_vector) return uint1440_t;
subtype int1440_t is signed(1439 downto 0);
constant int1440_t_SLV_LEN : integer := 1440;
function int1440_t_to_slv(x : int1440_t) return std_logic_vector;
function slv_to_int1440_t(x : std_logic_vector) return int1440_t;
subtype uint1441_t is unsigned(1440 downto 0);
constant uint1441_t_SLV_LEN : integer := 1441;
function uint1441_t_to_slv(x : uint1441_t) return std_logic_vector;
function slv_to_uint1441_t(x : std_logic_vector) return uint1441_t;
subtype int1441_t is signed(1440 downto 0);
constant int1441_t_SLV_LEN : integer := 1441;
function int1441_t_to_slv(x : int1441_t) return std_logic_vector;
function slv_to_int1441_t(x : std_logic_vector) return int1441_t;
subtype uint1442_t is unsigned(1441 downto 0);
constant uint1442_t_SLV_LEN : integer := 1442;
function uint1442_t_to_slv(x : uint1442_t) return std_logic_vector;
function slv_to_uint1442_t(x : std_logic_vector) return uint1442_t;
subtype int1442_t is signed(1441 downto 0);
constant int1442_t_SLV_LEN : integer := 1442;
function int1442_t_to_slv(x : int1442_t) return std_logic_vector;
function slv_to_int1442_t(x : std_logic_vector) return int1442_t;
subtype uint1443_t is unsigned(1442 downto 0);
constant uint1443_t_SLV_LEN : integer := 1443;
function uint1443_t_to_slv(x : uint1443_t) return std_logic_vector;
function slv_to_uint1443_t(x : std_logic_vector) return uint1443_t;
subtype int1443_t is signed(1442 downto 0);
constant int1443_t_SLV_LEN : integer := 1443;
function int1443_t_to_slv(x : int1443_t) return std_logic_vector;
function slv_to_int1443_t(x : std_logic_vector) return int1443_t;
subtype uint1444_t is unsigned(1443 downto 0);
constant uint1444_t_SLV_LEN : integer := 1444;
function uint1444_t_to_slv(x : uint1444_t) return std_logic_vector;
function slv_to_uint1444_t(x : std_logic_vector) return uint1444_t;
subtype int1444_t is signed(1443 downto 0);
constant int1444_t_SLV_LEN : integer := 1444;
function int1444_t_to_slv(x : int1444_t) return std_logic_vector;
function slv_to_int1444_t(x : std_logic_vector) return int1444_t;
subtype uint1445_t is unsigned(1444 downto 0);
constant uint1445_t_SLV_LEN : integer := 1445;
function uint1445_t_to_slv(x : uint1445_t) return std_logic_vector;
function slv_to_uint1445_t(x : std_logic_vector) return uint1445_t;
subtype int1445_t is signed(1444 downto 0);
constant int1445_t_SLV_LEN : integer := 1445;
function int1445_t_to_slv(x : int1445_t) return std_logic_vector;
function slv_to_int1445_t(x : std_logic_vector) return int1445_t;
subtype uint1446_t is unsigned(1445 downto 0);
constant uint1446_t_SLV_LEN : integer := 1446;
function uint1446_t_to_slv(x : uint1446_t) return std_logic_vector;
function slv_to_uint1446_t(x : std_logic_vector) return uint1446_t;
subtype int1446_t is signed(1445 downto 0);
constant int1446_t_SLV_LEN : integer := 1446;
function int1446_t_to_slv(x : int1446_t) return std_logic_vector;
function slv_to_int1446_t(x : std_logic_vector) return int1446_t;
subtype uint1447_t is unsigned(1446 downto 0);
constant uint1447_t_SLV_LEN : integer := 1447;
function uint1447_t_to_slv(x : uint1447_t) return std_logic_vector;
function slv_to_uint1447_t(x : std_logic_vector) return uint1447_t;
subtype int1447_t is signed(1446 downto 0);
constant int1447_t_SLV_LEN : integer := 1447;
function int1447_t_to_slv(x : int1447_t) return std_logic_vector;
function slv_to_int1447_t(x : std_logic_vector) return int1447_t;
subtype uint1448_t is unsigned(1447 downto 0);
constant uint1448_t_SLV_LEN : integer := 1448;
function uint1448_t_to_slv(x : uint1448_t) return std_logic_vector;
function slv_to_uint1448_t(x : std_logic_vector) return uint1448_t;
subtype int1448_t is signed(1447 downto 0);
constant int1448_t_SLV_LEN : integer := 1448;
function int1448_t_to_slv(x : int1448_t) return std_logic_vector;
function slv_to_int1448_t(x : std_logic_vector) return int1448_t;
subtype uint1449_t is unsigned(1448 downto 0);
constant uint1449_t_SLV_LEN : integer := 1449;
function uint1449_t_to_slv(x : uint1449_t) return std_logic_vector;
function slv_to_uint1449_t(x : std_logic_vector) return uint1449_t;
subtype int1449_t is signed(1448 downto 0);
constant int1449_t_SLV_LEN : integer := 1449;
function int1449_t_to_slv(x : int1449_t) return std_logic_vector;
function slv_to_int1449_t(x : std_logic_vector) return int1449_t;
subtype uint1450_t is unsigned(1449 downto 0);
constant uint1450_t_SLV_LEN : integer := 1450;
function uint1450_t_to_slv(x : uint1450_t) return std_logic_vector;
function slv_to_uint1450_t(x : std_logic_vector) return uint1450_t;
subtype int1450_t is signed(1449 downto 0);
constant int1450_t_SLV_LEN : integer := 1450;
function int1450_t_to_slv(x : int1450_t) return std_logic_vector;
function slv_to_int1450_t(x : std_logic_vector) return int1450_t;
subtype uint1451_t is unsigned(1450 downto 0);
constant uint1451_t_SLV_LEN : integer := 1451;
function uint1451_t_to_slv(x : uint1451_t) return std_logic_vector;
function slv_to_uint1451_t(x : std_logic_vector) return uint1451_t;
subtype int1451_t is signed(1450 downto 0);
constant int1451_t_SLV_LEN : integer := 1451;
function int1451_t_to_slv(x : int1451_t) return std_logic_vector;
function slv_to_int1451_t(x : std_logic_vector) return int1451_t;
subtype uint1452_t is unsigned(1451 downto 0);
constant uint1452_t_SLV_LEN : integer := 1452;
function uint1452_t_to_slv(x : uint1452_t) return std_logic_vector;
function slv_to_uint1452_t(x : std_logic_vector) return uint1452_t;
subtype int1452_t is signed(1451 downto 0);
constant int1452_t_SLV_LEN : integer := 1452;
function int1452_t_to_slv(x : int1452_t) return std_logic_vector;
function slv_to_int1452_t(x : std_logic_vector) return int1452_t;
subtype uint1453_t is unsigned(1452 downto 0);
constant uint1453_t_SLV_LEN : integer := 1453;
function uint1453_t_to_slv(x : uint1453_t) return std_logic_vector;
function slv_to_uint1453_t(x : std_logic_vector) return uint1453_t;
subtype int1453_t is signed(1452 downto 0);
constant int1453_t_SLV_LEN : integer := 1453;
function int1453_t_to_slv(x : int1453_t) return std_logic_vector;
function slv_to_int1453_t(x : std_logic_vector) return int1453_t;
subtype uint1454_t is unsigned(1453 downto 0);
constant uint1454_t_SLV_LEN : integer := 1454;
function uint1454_t_to_slv(x : uint1454_t) return std_logic_vector;
function slv_to_uint1454_t(x : std_logic_vector) return uint1454_t;
subtype int1454_t is signed(1453 downto 0);
constant int1454_t_SLV_LEN : integer := 1454;
function int1454_t_to_slv(x : int1454_t) return std_logic_vector;
function slv_to_int1454_t(x : std_logic_vector) return int1454_t;
subtype uint1455_t is unsigned(1454 downto 0);
constant uint1455_t_SLV_LEN : integer := 1455;
function uint1455_t_to_slv(x : uint1455_t) return std_logic_vector;
function slv_to_uint1455_t(x : std_logic_vector) return uint1455_t;
subtype int1455_t is signed(1454 downto 0);
constant int1455_t_SLV_LEN : integer := 1455;
function int1455_t_to_slv(x : int1455_t) return std_logic_vector;
function slv_to_int1455_t(x : std_logic_vector) return int1455_t;
subtype uint1456_t is unsigned(1455 downto 0);
constant uint1456_t_SLV_LEN : integer := 1456;
function uint1456_t_to_slv(x : uint1456_t) return std_logic_vector;
function slv_to_uint1456_t(x : std_logic_vector) return uint1456_t;
subtype int1456_t is signed(1455 downto 0);
constant int1456_t_SLV_LEN : integer := 1456;
function int1456_t_to_slv(x : int1456_t) return std_logic_vector;
function slv_to_int1456_t(x : std_logic_vector) return int1456_t;
subtype uint1457_t is unsigned(1456 downto 0);
constant uint1457_t_SLV_LEN : integer := 1457;
function uint1457_t_to_slv(x : uint1457_t) return std_logic_vector;
function slv_to_uint1457_t(x : std_logic_vector) return uint1457_t;
subtype int1457_t is signed(1456 downto 0);
constant int1457_t_SLV_LEN : integer := 1457;
function int1457_t_to_slv(x : int1457_t) return std_logic_vector;
function slv_to_int1457_t(x : std_logic_vector) return int1457_t;
subtype uint1458_t is unsigned(1457 downto 0);
constant uint1458_t_SLV_LEN : integer := 1458;
function uint1458_t_to_slv(x : uint1458_t) return std_logic_vector;
function slv_to_uint1458_t(x : std_logic_vector) return uint1458_t;
subtype int1458_t is signed(1457 downto 0);
constant int1458_t_SLV_LEN : integer := 1458;
function int1458_t_to_slv(x : int1458_t) return std_logic_vector;
function slv_to_int1458_t(x : std_logic_vector) return int1458_t;
subtype uint1459_t is unsigned(1458 downto 0);
constant uint1459_t_SLV_LEN : integer := 1459;
function uint1459_t_to_slv(x : uint1459_t) return std_logic_vector;
function slv_to_uint1459_t(x : std_logic_vector) return uint1459_t;
subtype int1459_t is signed(1458 downto 0);
constant int1459_t_SLV_LEN : integer := 1459;
function int1459_t_to_slv(x : int1459_t) return std_logic_vector;
function slv_to_int1459_t(x : std_logic_vector) return int1459_t;
subtype uint1460_t is unsigned(1459 downto 0);
constant uint1460_t_SLV_LEN : integer := 1460;
function uint1460_t_to_slv(x : uint1460_t) return std_logic_vector;
function slv_to_uint1460_t(x : std_logic_vector) return uint1460_t;
subtype int1460_t is signed(1459 downto 0);
constant int1460_t_SLV_LEN : integer := 1460;
function int1460_t_to_slv(x : int1460_t) return std_logic_vector;
function slv_to_int1460_t(x : std_logic_vector) return int1460_t;
subtype uint1461_t is unsigned(1460 downto 0);
constant uint1461_t_SLV_LEN : integer := 1461;
function uint1461_t_to_slv(x : uint1461_t) return std_logic_vector;
function slv_to_uint1461_t(x : std_logic_vector) return uint1461_t;
subtype int1461_t is signed(1460 downto 0);
constant int1461_t_SLV_LEN : integer := 1461;
function int1461_t_to_slv(x : int1461_t) return std_logic_vector;
function slv_to_int1461_t(x : std_logic_vector) return int1461_t;
subtype uint1462_t is unsigned(1461 downto 0);
constant uint1462_t_SLV_LEN : integer := 1462;
function uint1462_t_to_slv(x : uint1462_t) return std_logic_vector;
function slv_to_uint1462_t(x : std_logic_vector) return uint1462_t;
subtype int1462_t is signed(1461 downto 0);
constant int1462_t_SLV_LEN : integer := 1462;
function int1462_t_to_slv(x : int1462_t) return std_logic_vector;
function slv_to_int1462_t(x : std_logic_vector) return int1462_t;
subtype uint1463_t is unsigned(1462 downto 0);
constant uint1463_t_SLV_LEN : integer := 1463;
function uint1463_t_to_slv(x : uint1463_t) return std_logic_vector;
function slv_to_uint1463_t(x : std_logic_vector) return uint1463_t;
subtype int1463_t is signed(1462 downto 0);
constant int1463_t_SLV_LEN : integer := 1463;
function int1463_t_to_slv(x : int1463_t) return std_logic_vector;
function slv_to_int1463_t(x : std_logic_vector) return int1463_t;
subtype uint1464_t is unsigned(1463 downto 0);
constant uint1464_t_SLV_LEN : integer := 1464;
function uint1464_t_to_slv(x : uint1464_t) return std_logic_vector;
function slv_to_uint1464_t(x : std_logic_vector) return uint1464_t;
subtype int1464_t is signed(1463 downto 0);
constant int1464_t_SLV_LEN : integer := 1464;
function int1464_t_to_slv(x : int1464_t) return std_logic_vector;
function slv_to_int1464_t(x : std_logic_vector) return int1464_t;
subtype uint1465_t is unsigned(1464 downto 0);
constant uint1465_t_SLV_LEN : integer := 1465;
function uint1465_t_to_slv(x : uint1465_t) return std_logic_vector;
function slv_to_uint1465_t(x : std_logic_vector) return uint1465_t;
subtype int1465_t is signed(1464 downto 0);
constant int1465_t_SLV_LEN : integer := 1465;
function int1465_t_to_slv(x : int1465_t) return std_logic_vector;
function slv_to_int1465_t(x : std_logic_vector) return int1465_t;
subtype uint1466_t is unsigned(1465 downto 0);
constant uint1466_t_SLV_LEN : integer := 1466;
function uint1466_t_to_slv(x : uint1466_t) return std_logic_vector;
function slv_to_uint1466_t(x : std_logic_vector) return uint1466_t;
subtype int1466_t is signed(1465 downto 0);
constant int1466_t_SLV_LEN : integer := 1466;
function int1466_t_to_slv(x : int1466_t) return std_logic_vector;
function slv_to_int1466_t(x : std_logic_vector) return int1466_t;
subtype uint1467_t is unsigned(1466 downto 0);
constant uint1467_t_SLV_LEN : integer := 1467;
function uint1467_t_to_slv(x : uint1467_t) return std_logic_vector;
function slv_to_uint1467_t(x : std_logic_vector) return uint1467_t;
subtype int1467_t is signed(1466 downto 0);
constant int1467_t_SLV_LEN : integer := 1467;
function int1467_t_to_slv(x : int1467_t) return std_logic_vector;
function slv_to_int1467_t(x : std_logic_vector) return int1467_t;
subtype uint1468_t is unsigned(1467 downto 0);
constant uint1468_t_SLV_LEN : integer := 1468;
function uint1468_t_to_slv(x : uint1468_t) return std_logic_vector;
function slv_to_uint1468_t(x : std_logic_vector) return uint1468_t;
subtype int1468_t is signed(1467 downto 0);
constant int1468_t_SLV_LEN : integer := 1468;
function int1468_t_to_slv(x : int1468_t) return std_logic_vector;
function slv_to_int1468_t(x : std_logic_vector) return int1468_t;
subtype uint1469_t is unsigned(1468 downto 0);
constant uint1469_t_SLV_LEN : integer := 1469;
function uint1469_t_to_slv(x : uint1469_t) return std_logic_vector;
function slv_to_uint1469_t(x : std_logic_vector) return uint1469_t;
subtype int1469_t is signed(1468 downto 0);
constant int1469_t_SLV_LEN : integer := 1469;
function int1469_t_to_slv(x : int1469_t) return std_logic_vector;
function slv_to_int1469_t(x : std_logic_vector) return int1469_t;
subtype uint1470_t is unsigned(1469 downto 0);
constant uint1470_t_SLV_LEN : integer := 1470;
function uint1470_t_to_slv(x : uint1470_t) return std_logic_vector;
function slv_to_uint1470_t(x : std_logic_vector) return uint1470_t;
subtype int1470_t is signed(1469 downto 0);
constant int1470_t_SLV_LEN : integer := 1470;
function int1470_t_to_slv(x : int1470_t) return std_logic_vector;
function slv_to_int1470_t(x : std_logic_vector) return int1470_t;
subtype uint1471_t is unsigned(1470 downto 0);
constant uint1471_t_SLV_LEN : integer := 1471;
function uint1471_t_to_slv(x : uint1471_t) return std_logic_vector;
function slv_to_uint1471_t(x : std_logic_vector) return uint1471_t;
subtype int1471_t is signed(1470 downto 0);
constant int1471_t_SLV_LEN : integer := 1471;
function int1471_t_to_slv(x : int1471_t) return std_logic_vector;
function slv_to_int1471_t(x : std_logic_vector) return int1471_t;
subtype uint1472_t is unsigned(1471 downto 0);
constant uint1472_t_SLV_LEN : integer := 1472;
function uint1472_t_to_slv(x : uint1472_t) return std_logic_vector;
function slv_to_uint1472_t(x : std_logic_vector) return uint1472_t;
subtype int1472_t is signed(1471 downto 0);
constant int1472_t_SLV_LEN : integer := 1472;
function int1472_t_to_slv(x : int1472_t) return std_logic_vector;
function slv_to_int1472_t(x : std_logic_vector) return int1472_t;
subtype uint1473_t is unsigned(1472 downto 0);
constant uint1473_t_SLV_LEN : integer := 1473;
function uint1473_t_to_slv(x : uint1473_t) return std_logic_vector;
function slv_to_uint1473_t(x : std_logic_vector) return uint1473_t;
subtype int1473_t is signed(1472 downto 0);
constant int1473_t_SLV_LEN : integer := 1473;
function int1473_t_to_slv(x : int1473_t) return std_logic_vector;
function slv_to_int1473_t(x : std_logic_vector) return int1473_t;
subtype uint1474_t is unsigned(1473 downto 0);
constant uint1474_t_SLV_LEN : integer := 1474;
function uint1474_t_to_slv(x : uint1474_t) return std_logic_vector;
function slv_to_uint1474_t(x : std_logic_vector) return uint1474_t;
subtype int1474_t is signed(1473 downto 0);
constant int1474_t_SLV_LEN : integer := 1474;
function int1474_t_to_slv(x : int1474_t) return std_logic_vector;
function slv_to_int1474_t(x : std_logic_vector) return int1474_t;
subtype uint1475_t is unsigned(1474 downto 0);
constant uint1475_t_SLV_LEN : integer := 1475;
function uint1475_t_to_slv(x : uint1475_t) return std_logic_vector;
function slv_to_uint1475_t(x : std_logic_vector) return uint1475_t;
subtype int1475_t is signed(1474 downto 0);
constant int1475_t_SLV_LEN : integer := 1475;
function int1475_t_to_slv(x : int1475_t) return std_logic_vector;
function slv_to_int1475_t(x : std_logic_vector) return int1475_t;
subtype uint1476_t is unsigned(1475 downto 0);
constant uint1476_t_SLV_LEN : integer := 1476;
function uint1476_t_to_slv(x : uint1476_t) return std_logic_vector;
function slv_to_uint1476_t(x : std_logic_vector) return uint1476_t;
subtype int1476_t is signed(1475 downto 0);
constant int1476_t_SLV_LEN : integer := 1476;
function int1476_t_to_slv(x : int1476_t) return std_logic_vector;
function slv_to_int1476_t(x : std_logic_vector) return int1476_t;
subtype uint1477_t is unsigned(1476 downto 0);
constant uint1477_t_SLV_LEN : integer := 1477;
function uint1477_t_to_slv(x : uint1477_t) return std_logic_vector;
function slv_to_uint1477_t(x : std_logic_vector) return uint1477_t;
subtype int1477_t is signed(1476 downto 0);
constant int1477_t_SLV_LEN : integer := 1477;
function int1477_t_to_slv(x : int1477_t) return std_logic_vector;
function slv_to_int1477_t(x : std_logic_vector) return int1477_t;
subtype uint1478_t is unsigned(1477 downto 0);
constant uint1478_t_SLV_LEN : integer := 1478;
function uint1478_t_to_slv(x : uint1478_t) return std_logic_vector;
function slv_to_uint1478_t(x : std_logic_vector) return uint1478_t;
subtype int1478_t is signed(1477 downto 0);
constant int1478_t_SLV_LEN : integer := 1478;
function int1478_t_to_slv(x : int1478_t) return std_logic_vector;
function slv_to_int1478_t(x : std_logic_vector) return int1478_t;
subtype uint1479_t is unsigned(1478 downto 0);
constant uint1479_t_SLV_LEN : integer := 1479;
function uint1479_t_to_slv(x : uint1479_t) return std_logic_vector;
function slv_to_uint1479_t(x : std_logic_vector) return uint1479_t;
subtype int1479_t is signed(1478 downto 0);
constant int1479_t_SLV_LEN : integer := 1479;
function int1479_t_to_slv(x : int1479_t) return std_logic_vector;
function slv_to_int1479_t(x : std_logic_vector) return int1479_t;
subtype uint1480_t is unsigned(1479 downto 0);
constant uint1480_t_SLV_LEN : integer := 1480;
function uint1480_t_to_slv(x : uint1480_t) return std_logic_vector;
function slv_to_uint1480_t(x : std_logic_vector) return uint1480_t;
subtype int1480_t is signed(1479 downto 0);
constant int1480_t_SLV_LEN : integer := 1480;
function int1480_t_to_slv(x : int1480_t) return std_logic_vector;
function slv_to_int1480_t(x : std_logic_vector) return int1480_t;
subtype uint1481_t is unsigned(1480 downto 0);
constant uint1481_t_SLV_LEN : integer := 1481;
function uint1481_t_to_slv(x : uint1481_t) return std_logic_vector;
function slv_to_uint1481_t(x : std_logic_vector) return uint1481_t;
subtype int1481_t is signed(1480 downto 0);
constant int1481_t_SLV_LEN : integer := 1481;
function int1481_t_to_slv(x : int1481_t) return std_logic_vector;
function slv_to_int1481_t(x : std_logic_vector) return int1481_t;
subtype uint1482_t is unsigned(1481 downto 0);
constant uint1482_t_SLV_LEN : integer := 1482;
function uint1482_t_to_slv(x : uint1482_t) return std_logic_vector;
function slv_to_uint1482_t(x : std_logic_vector) return uint1482_t;
subtype int1482_t is signed(1481 downto 0);
constant int1482_t_SLV_LEN : integer := 1482;
function int1482_t_to_slv(x : int1482_t) return std_logic_vector;
function slv_to_int1482_t(x : std_logic_vector) return int1482_t;
subtype uint1483_t is unsigned(1482 downto 0);
constant uint1483_t_SLV_LEN : integer := 1483;
function uint1483_t_to_slv(x : uint1483_t) return std_logic_vector;
function slv_to_uint1483_t(x : std_logic_vector) return uint1483_t;
subtype int1483_t is signed(1482 downto 0);
constant int1483_t_SLV_LEN : integer := 1483;
function int1483_t_to_slv(x : int1483_t) return std_logic_vector;
function slv_to_int1483_t(x : std_logic_vector) return int1483_t;
subtype uint1484_t is unsigned(1483 downto 0);
constant uint1484_t_SLV_LEN : integer := 1484;
function uint1484_t_to_slv(x : uint1484_t) return std_logic_vector;
function slv_to_uint1484_t(x : std_logic_vector) return uint1484_t;
subtype int1484_t is signed(1483 downto 0);
constant int1484_t_SLV_LEN : integer := 1484;
function int1484_t_to_slv(x : int1484_t) return std_logic_vector;
function slv_to_int1484_t(x : std_logic_vector) return int1484_t;
subtype uint1485_t is unsigned(1484 downto 0);
constant uint1485_t_SLV_LEN : integer := 1485;
function uint1485_t_to_slv(x : uint1485_t) return std_logic_vector;
function slv_to_uint1485_t(x : std_logic_vector) return uint1485_t;
subtype int1485_t is signed(1484 downto 0);
constant int1485_t_SLV_LEN : integer := 1485;
function int1485_t_to_slv(x : int1485_t) return std_logic_vector;
function slv_to_int1485_t(x : std_logic_vector) return int1485_t;
subtype uint1486_t is unsigned(1485 downto 0);
constant uint1486_t_SLV_LEN : integer := 1486;
function uint1486_t_to_slv(x : uint1486_t) return std_logic_vector;
function slv_to_uint1486_t(x : std_logic_vector) return uint1486_t;
subtype int1486_t is signed(1485 downto 0);
constant int1486_t_SLV_LEN : integer := 1486;
function int1486_t_to_slv(x : int1486_t) return std_logic_vector;
function slv_to_int1486_t(x : std_logic_vector) return int1486_t;
subtype uint1487_t is unsigned(1486 downto 0);
constant uint1487_t_SLV_LEN : integer := 1487;
function uint1487_t_to_slv(x : uint1487_t) return std_logic_vector;
function slv_to_uint1487_t(x : std_logic_vector) return uint1487_t;
subtype int1487_t is signed(1486 downto 0);
constant int1487_t_SLV_LEN : integer := 1487;
function int1487_t_to_slv(x : int1487_t) return std_logic_vector;
function slv_to_int1487_t(x : std_logic_vector) return int1487_t;
subtype uint1488_t is unsigned(1487 downto 0);
constant uint1488_t_SLV_LEN : integer := 1488;
function uint1488_t_to_slv(x : uint1488_t) return std_logic_vector;
function slv_to_uint1488_t(x : std_logic_vector) return uint1488_t;
subtype int1488_t is signed(1487 downto 0);
constant int1488_t_SLV_LEN : integer := 1488;
function int1488_t_to_slv(x : int1488_t) return std_logic_vector;
function slv_to_int1488_t(x : std_logic_vector) return int1488_t;
subtype uint1489_t is unsigned(1488 downto 0);
constant uint1489_t_SLV_LEN : integer := 1489;
function uint1489_t_to_slv(x : uint1489_t) return std_logic_vector;
function slv_to_uint1489_t(x : std_logic_vector) return uint1489_t;
subtype int1489_t is signed(1488 downto 0);
constant int1489_t_SLV_LEN : integer := 1489;
function int1489_t_to_slv(x : int1489_t) return std_logic_vector;
function slv_to_int1489_t(x : std_logic_vector) return int1489_t;
subtype uint1490_t is unsigned(1489 downto 0);
constant uint1490_t_SLV_LEN : integer := 1490;
function uint1490_t_to_slv(x : uint1490_t) return std_logic_vector;
function slv_to_uint1490_t(x : std_logic_vector) return uint1490_t;
subtype int1490_t is signed(1489 downto 0);
constant int1490_t_SLV_LEN : integer := 1490;
function int1490_t_to_slv(x : int1490_t) return std_logic_vector;
function slv_to_int1490_t(x : std_logic_vector) return int1490_t;
subtype uint1491_t is unsigned(1490 downto 0);
constant uint1491_t_SLV_LEN : integer := 1491;
function uint1491_t_to_slv(x : uint1491_t) return std_logic_vector;
function slv_to_uint1491_t(x : std_logic_vector) return uint1491_t;
subtype int1491_t is signed(1490 downto 0);
constant int1491_t_SLV_LEN : integer := 1491;
function int1491_t_to_slv(x : int1491_t) return std_logic_vector;
function slv_to_int1491_t(x : std_logic_vector) return int1491_t;
subtype uint1492_t is unsigned(1491 downto 0);
constant uint1492_t_SLV_LEN : integer := 1492;
function uint1492_t_to_slv(x : uint1492_t) return std_logic_vector;
function slv_to_uint1492_t(x : std_logic_vector) return uint1492_t;
subtype int1492_t is signed(1491 downto 0);
constant int1492_t_SLV_LEN : integer := 1492;
function int1492_t_to_slv(x : int1492_t) return std_logic_vector;
function slv_to_int1492_t(x : std_logic_vector) return int1492_t;
subtype uint1493_t is unsigned(1492 downto 0);
constant uint1493_t_SLV_LEN : integer := 1493;
function uint1493_t_to_slv(x : uint1493_t) return std_logic_vector;
function slv_to_uint1493_t(x : std_logic_vector) return uint1493_t;
subtype int1493_t is signed(1492 downto 0);
constant int1493_t_SLV_LEN : integer := 1493;
function int1493_t_to_slv(x : int1493_t) return std_logic_vector;
function slv_to_int1493_t(x : std_logic_vector) return int1493_t;
subtype uint1494_t is unsigned(1493 downto 0);
constant uint1494_t_SLV_LEN : integer := 1494;
function uint1494_t_to_slv(x : uint1494_t) return std_logic_vector;
function slv_to_uint1494_t(x : std_logic_vector) return uint1494_t;
subtype int1494_t is signed(1493 downto 0);
constant int1494_t_SLV_LEN : integer := 1494;
function int1494_t_to_slv(x : int1494_t) return std_logic_vector;
function slv_to_int1494_t(x : std_logic_vector) return int1494_t;
subtype uint1495_t is unsigned(1494 downto 0);
constant uint1495_t_SLV_LEN : integer := 1495;
function uint1495_t_to_slv(x : uint1495_t) return std_logic_vector;
function slv_to_uint1495_t(x : std_logic_vector) return uint1495_t;
subtype int1495_t is signed(1494 downto 0);
constant int1495_t_SLV_LEN : integer := 1495;
function int1495_t_to_slv(x : int1495_t) return std_logic_vector;
function slv_to_int1495_t(x : std_logic_vector) return int1495_t;
subtype uint1496_t is unsigned(1495 downto 0);
constant uint1496_t_SLV_LEN : integer := 1496;
function uint1496_t_to_slv(x : uint1496_t) return std_logic_vector;
function slv_to_uint1496_t(x : std_logic_vector) return uint1496_t;
subtype int1496_t is signed(1495 downto 0);
constant int1496_t_SLV_LEN : integer := 1496;
function int1496_t_to_slv(x : int1496_t) return std_logic_vector;
function slv_to_int1496_t(x : std_logic_vector) return int1496_t;
subtype uint1497_t is unsigned(1496 downto 0);
constant uint1497_t_SLV_LEN : integer := 1497;
function uint1497_t_to_slv(x : uint1497_t) return std_logic_vector;
function slv_to_uint1497_t(x : std_logic_vector) return uint1497_t;
subtype int1497_t is signed(1496 downto 0);
constant int1497_t_SLV_LEN : integer := 1497;
function int1497_t_to_slv(x : int1497_t) return std_logic_vector;
function slv_to_int1497_t(x : std_logic_vector) return int1497_t;
subtype uint1498_t is unsigned(1497 downto 0);
constant uint1498_t_SLV_LEN : integer := 1498;
function uint1498_t_to_slv(x : uint1498_t) return std_logic_vector;
function slv_to_uint1498_t(x : std_logic_vector) return uint1498_t;
subtype int1498_t is signed(1497 downto 0);
constant int1498_t_SLV_LEN : integer := 1498;
function int1498_t_to_slv(x : int1498_t) return std_logic_vector;
function slv_to_int1498_t(x : std_logic_vector) return int1498_t;
subtype uint1499_t is unsigned(1498 downto 0);
constant uint1499_t_SLV_LEN : integer := 1499;
function uint1499_t_to_slv(x : uint1499_t) return std_logic_vector;
function slv_to_uint1499_t(x : std_logic_vector) return uint1499_t;
subtype int1499_t is signed(1498 downto 0);
constant int1499_t_SLV_LEN : integer := 1499;
function int1499_t_to_slv(x : int1499_t) return std_logic_vector;
function slv_to_int1499_t(x : std_logic_vector) return int1499_t;
subtype uint1500_t is unsigned(1499 downto 0);
constant uint1500_t_SLV_LEN : integer := 1500;
function uint1500_t_to_slv(x : uint1500_t) return std_logic_vector;
function slv_to_uint1500_t(x : std_logic_vector) return uint1500_t;
subtype int1500_t is signed(1499 downto 0);
constant int1500_t_SLV_LEN : integer := 1500;
function int1500_t_to_slv(x : int1500_t) return std_logic_vector;
function slv_to_int1500_t(x : std_logic_vector) return int1500_t;
subtype uint1501_t is unsigned(1500 downto 0);
constant uint1501_t_SLV_LEN : integer := 1501;
function uint1501_t_to_slv(x : uint1501_t) return std_logic_vector;
function slv_to_uint1501_t(x : std_logic_vector) return uint1501_t;
subtype int1501_t is signed(1500 downto 0);
constant int1501_t_SLV_LEN : integer := 1501;
function int1501_t_to_slv(x : int1501_t) return std_logic_vector;
function slv_to_int1501_t(x : std_logic_vector) return int1501_t;
subtype uint1502_t is unsigned(1501 downto 0);
constant uint1502_t_SLV_LEN : integer := 1502;
function uint1502_t_to_slv(x : uint1502_t) return std_logic_vector;
function slv_to_uint1502_t(x : std_logic_vector) return uint1502_t;
subtype int1502_t is signed(1501 downto 0);
constant int1502_t_SLV_LEN : integer := 1502;
function int1502_t_to_slv(x : int1502_t) return std_logic_vector;
function slv_to_int1502_t(x : std_logic_vector) return int1502_t;
subtype uint1503_t is unsigned(1502 downto 0);
constant uint1503_t_SLV_LEN : integer := 1503;
function uint1503_t_to_slv(x : uint1503_t) return std_logic_vector;
function slv_to_uint1503_t(x : std_logic_vector) return uint1503_t;
subtype int1503_t is signed(1502 downto 0);
constant int1503_t_SLV_LEN : integer := 1503;
function int1503_t_to_slv(x : int1503_t) return std_logic_vector;
function slv_to_int1503_t(x : std_logic_vector) return int1503_t;
subtype uint1504_t is unsigned(1503 downto 0);
constant uint1504_t_SLV_LEN : integer := 1504;
function uint1504_t_to_slv(x : uint1504_t) return std_logic_vector;
function slv_to_uint1504_t(x : std_logic_vector) return uint1504_t;
subtype int1504_t is signed(1503 downto 0);
constant int1504_t_SLV_LEN : integer := 1504;
function int1504_t_to_slv(x : int1504_t) return std_logic_vector;
function slv_to_int1504_t(x : std_logic_vector) return int1504_t;
subtype uint1505_t is unsigned(1504 downto 0);
constant uint1505_t_SLV_LEN : integer := 1505;
function uint1505_t_to_slv(x : uint1505_t) return std_logic_vector;
function slv_to_uint1505_t(x : std_logic_vector) return uint1505_t;
subtype int1505_t is signed(1504 downto 0);
constant int1505_t_SLV_LEN : integer := 1505;
function int1505_t_to_slv(x : int1505_t) return std_logic_vector;
function slv_to_int1505_t(x : std_logic_vector) return int1505_t;
subtype uint1506_t is unsigned(1505 downto 0);
constant uint1506_t_SLV_LEN : integer := 1506;
function uint1506_t_to_slv(x : uint1506_t) return std_logic_vector;
function slv_to_uint1506_t(x : std_logic_vector) return uint1506_t;
subtype int1506_t is signed(1505 downto 0);
constant int1506_t_SLV_LEN : integer := 1506;
function int1506_t_to_slv(x : int1506_t) return std_logic_vector;
function slv_to_int1506_t(x : std_logic_vector) return int1506_t;
subtype uint1507_t is unsigned(1506 downto 0);
constant uint1507_t_SLV_LEN : integer := 1507;
function uint1507_t_to_slv(x : uint1507_t) return std_logic_vector;
function slv_to_uint1507_t(x : std_logic_vector) return uint1507_t;
subtype int1507_t is signed(1506 downto 0);
constant int1507_t_SLV_LEN : integer := 1507;
function int1507_t_to_slv(x : int1507_t) return std_logic_vector;
function slv_to_int1507_t(x : std_logic_vector) return int1507_t;
subtype uint1508_t is unsigned(1507 downto 0);
constant uint1508_t_SLV_LEN : integer := 1508;
function uint1508_t_to_slv(x : uint1508_t) return std_logic_vector;
function slv_to_uint1508_t(x : std_logic_vector) return uint1508_t;
subtype int1508_t is signed(1507 downto 0);
constant int1508_t_SLV_LEN : integer := 1508;
function int1508_t_to_slv(x : int1508_t) return std_logic_vector;
function slv_to_int1508_t(x : std_logic_vector) return int1508_t;
subtype uint1509_t is unsigned(1508 downto 0);
constant uint1509_t_SLV_LEN : integer := 1509;
function uint1509_t_to_slv(x : uint1509_t) return std_logic_vector;
function slv_to_uint1509_t(x : std_logic_vector) return uint1509_t;
subtype int1509_t is signed(1508 downto 0);
constant int1509_t_SLV_LEN : integer := 1509;
function int1509_t_to_slv(x : int1509_t) return std_logic_vector;
function slv_to_int1509_t(x : std_logic_vector) return int1509_t;
subtype uint1510_t is unsigned(1509 downto 0);
constant uint1510_t_SLV_LEN : integer := 1510;
function uint1510_t_to_slv(x : uint1510_t) return std_logic_vector;
function slv_to_uint1510_t(x : std_logic_vector) return uint1510_t;
subtype int1510_t is signed(1509 downto 0);
constant int1510_t_SLV_LEN : integer := 1510;
function int1510_t_to_slv(x : int1510_t) return std_logic_vector;
function slv_to_int1510_t(x : std_logic_vector) return int1510_t;
subtype uint1511_t is unsigned(1510 downto 0);
constant uint1511_t_SLV_LEN : integer := 1511;
function uint1511_t_to_slv(x : uint1511_t) return std_logic_vector;
function slv_to_uint1511_t(x : std_logic_vector) return uint1511_t;
subtype int1511_t is signed(1510 downto 0);
constant int1511_t_SLV_LEN : integer := 1511;
function int1511_t_to_slv(x : int1511_t) return std_logic_vector;
function slv_to_int1511_t(x : std_logic_vector) return int1511_t;
subtype uint1512_t is unsigned(1511 downto 0);
constant uint1512_t_SLV_LEN : integer := 1512;
function uint1512_t_to_slv(x : uint1512_t) return std_logic_vector;
function slv_to_uint1512_t(x : std_logic_vector) return uint1512_t;
subtype int1512_t is signed(1511 downto 0);
constant int1512_t_SLV_LEN : integer := 1512;
function int1512_t_to_slv(x : int1512_t) return std_logic_vector;
function slv_to_int1512_t(x : std_logic_vector) return int1512_t;
subtype uint1513_t is unsigned(1512 downto 0);
constant uint1513_t_SLV_LEN : integer := 1513;
function uint1513_t_to_slv(x : uint1513_t) return std_logic_vector;
function slv_to_uint1513_t(x : std_logic_vector) return uint1513_t;
subtype int1513_t is signed(1512 downto 0);
constant int1513_t_SLV_LEN : integer := 1513;
function int1513_t_to_slv(x : int1513_t) return std_logic_vector;
function slv_to_int1513_t(x : std_logic_vector) return int1513_t;
subtype uint1514_t is unsigned(1513 downto 0);
constant uint1514_t_SLV_LEN : integer := 1514;
function uint1514_t_to_slv(x : uint1514_t) return std_logic_vector;
function slv_to_uint1514_t(x : std_logic_vector) return uint1514_t;
subtype int1514_t is signed(1513 downto 0);
constant int1514_t_SLV_LEN : integer := 1514;
function int1514_t_to_slv(x : int1514_t) return std_logic_vector;
function slv_to_int1514_t(x : std_logic_vector) return int1514_t;
subtype uint1515_t is unsigned(1514 downto 0);
constant uint1515_t_SLV_LEN : integer := 1515;
function uint1515_t_to_slv(x : uint1515_t) return std_logic_vector;
function slv_to_uint1515_t(x : std_logic_vector) return uint1515_t;
subtype int1515_t is signed(1514 downto 0);
constant int1515_t_SLV_LEN : integer := 1515;
function int1515_t_to_slv(x : int1515_t) return std_logic_vector;
function slv_to_int1515_t(x : std_logic_vector) return int1515_t;
subtype uint1516_t is unsigned(1515 downto 0);
constant uint1516_t_SLV_LEN : integer := 1516;
function uint1516_t_to_slv(x : uint1516_t) return std_logic_vector;
function slv_to_uint1516_t(x : std_logic_vector) return uint1516_t;
subtype int1516_t is signed(1515 downto 0);
constant int1516_t_SLV_LEN : integer := 1516;
function int1516_t_to_slv(x : int1516_t) return std_logic_vector;
function slv_to_int1516_t(x : std_logic_vector) return int1516_t;
subtype uint1517_t is unsigned(1516 downto 0);
constant uint1517_t_SLV_LEN : integer := 1517;
function uint1517_t_to_slv(x : uint1517_t) return std_logic_vector;
function slv_to_uint1517_t(x : std_logic_vector) return uint1517_t;
subtype int1517_t is signed(1516 downto 0);
constant int1517_t_SLV_LEN : integer := 1517;
function int1517_t_to_slv(x : int1517_t) return std_logic_vector;
function slv_to_int1517_t(x : std_logic_vector) return int1517_t;
subtype uint1518_t is unsigned(1517 downto 0);
constant uint1518_t_SLV_LEN : integer := 1518;
function uint1518_t_to_slv(x : uint1518_t) return std_logic_vector;
function slv_to_uint1518_t(x : std_logic_vector) return uint1518_t;
subtype int1518_t is signed(1517 downto 0);
constant int1518_t_SLV_LEN : integer := 1518;
function int1518_t_to_slv(x : int1518_t) return std_logic_vector;
function slv_to_int1518_t(x : std_logic_vector) return int1518_t;
subtype uint1519_t is unsigned(1518 downto 0);
constant uint1519_t_SLV_LEN : integer := 1519;
function uint1519_t_to_slv(x : uint1519_t) return std_logic_vector;
function slv_to_uint1519_t(x : std_logic_vector) return uint1519_t;
subtype int1519_t is signed(1518 downto 0);
constant int1519_t_SLV_LEN : integer := 1519;
function int1519_t_to_slv(x : int1519_t) return std_logic_vector;
function slv_to_int1519_t(x : std_logic_vector) return int1519_t;
subtype uint1520_t is unsigned(1519 downto 0);
constant uint1520_t_SLV_LEN : integer := 1520;
function uint1520_t_to_slv(x : uint1520_t) return std_logic_vector;
function slv_to_uint1520_t(x : std_logic_vector) return uint1520_t;
subtype int1520_t is signed(1519 downto 0);
constant int1520_t_SLV_LEN : integer := 1520;
function int1520_t_to_slv(x : int1520_t) return std_logic_vector;
function slv_to_int1520_t(x : std_logic_vector) return int1520_t;
subtype uint1521_t is unsigned(1520 downto 0);
constant uint1521_t_SLV_LEN : integer := 1521;
function uint1521_t_to_slv(x : uint1521_t) return std_logic_vector;
function slv_to_uint1521_t(x : std_logic_vector) return uint1521_t;
subtype int1521_t is signed(1520 downto 0);
constant int1521_t_SLV_LEN : integer := 1521;
function int1521_t_to_slv(x : int1521_t) return std_logic_vector;
function slv_to_int1521_t(x : std_logic_vector) return int1521_t;
subtype uint1522_t is unsigned(1521 downto 0);
constant uint1522_t_SLV_LEN : integer := 1522;
function uint1522_t_to_slv(x : uint1522_t) return std_logic_vector;
function slv_to_uint1522_t(x : std_logic_vector) return uint1522_t;
subtype int1522_t is signed(1521 downto 0);
constant int1522_t_SLV_LEN : integer := 1522;
function int1522_t_to_slv(x : int1522_t) return std_logic_vector;
function slv_to_int1522_t(x : std_logic_vector) return int1522_t;
subtype uint1523_t is unsigned(1522 downto 0);
constant uint1523_t_SLV_LEN : integer := 1523;
function uint1523_t_to_slv(x : uint1523_t) return std_logic_vector;
function slv_to_uint1523_t(x : std_logic_vector) return uint1523_t;
subtype int1523_t is signed(1522 downto 0);
constant int1523_t_SLV_LEN : integer := 1523;
function int1523_t_to_slv(x : int1523_t) return std_logic_vector;
function slv_to_int1523_t(x : std_logic_vector) return int1523_t;
subtype uint1524_t is unsigned(1523 downto 0);
constant uint1524_t_SLV_LEN : integer := 1524;
function uint1524_t_to_slv(x : uint1524_t) return std_logic_vector;
function slv_to_uint1524_t(x : std_logic_vector) return uint1524_t;
subtype int1524_t is signed(1523 downto 0);
constant int1524_t_SLV_LEN : integer := 1524;
function int1524_t_to_slv(x : int1524_t) return std_logic_vector;
function slv_to_int1524_t(x : std_logic_vector) return int1524_t;
subtype uint1525_t is unsigned(1524 downto 0);
constant uint1525_t_SLV_LEN : integer := 1525;
function uint1525_t_to_slv(x : uint1525_t) return std_logic_vector;
function slv_to_uint1525_t(x : std_logic_vector) return uint1525_t;
subtype int1525_t is signed(1524 downto 0);
constant int1525_t_SLV_LEN : integer := 1525;
function int1525_t_to_slv(x : int1525_t) return std_logic_vector;
function slv_to_int1525_t(x : std_logic_vector) return int1525_t;
subtype uint1526_t is unsigned(1525 downto 0);
constant uint1526_t_SLV_LEN : integer := 1526;
function uint1526_t_to_slv(x : uint1526_t) return std_logic_vector;
function slv_to_uint1526_t(x : std_logic_vector) return uint1526_t;
subtype int1526_t is signed(1525 downto 0);
constant int1526_t_SLV_LEN : integer := 1526;
function int1526_t_to_slv(x : int1526_t) return std_logic_vector;
function slv_to_int1526_t(x : std_logic_vector) return int1526_t;
subtype uint1527_t is unsigned(1526 downto 0);
constant uint1527_t_SLV_LEN : integer := 1527;
function uint1527_t_to_slv(x : uint1527_t) return std_logic_vector;
function slv_to_uint1527_t(x : std_logic_vector) return uint1527_t;
subtype int1527_t is signed(1526 downto 0);
constant int1527_t_SLV_LEN : integer := 1527;
function int1527_t_to_slv(x : int1527_t) return std_logic_vector;
function slv_to_int1527_t(x : std_logic_vector) return int1527_t;
subtype uint1528_t is unsigned(1527 downto 0);
constant uint1528_t_SLV_LEN : integer := 1528;
function uint1528_t_to_slv(x : uint1528_t) return std_logic_vector;
function slv_to_uint1528_t(x : std_logic_vector) return uint1528_t;
subtype int1528_t is signed(1527 downto 0);
constant int1528_t_SLV_LEN : integer := 1528;
function int1528_t_to_slv(x : int1528_t) return std_logic_vector;
function slv_to_int1528_t(x : std_logic_vector) return int1528_t;
subtype uint1529_t is unsigned(1528 downto 0);
constant uint1529_t_SLV_LEN : integer := 1529;
function uint1529_t_to_slv(x : uint1529_t) return std_logic_vector;
function slv_to_uint1529_t(x : std_logic_vector) return uint1529_t;
subtype int1529_t is signed(1528 downto 0);
constant int1529_t_SLV_LEN : integer := 1529;
function int1529_t_to_slv(x : int1529_t) return std_logic_vector;
function slv_to_int1529_t(x : std_logic_vector) return int1529_t;
subtype uint1530_t is unsigned(1529 downto 0);
constant uint1530_t_SLV_LEN : integer := 1530;
function uint1530_t_to_slv(x : uint1530_t) return std_logic_vector;
function slv_to_uint1530_t(x : std_logic_vector) return uint1530_t;
subtype int1530_t is signed(1529 downto 0);
constant int1530_t_SLV_LEN : integer := 1530;
function int1530_t_to_slv(x : int1530_t) return std_logic_vector;
function slv_to_int1530_t(x : std_logic_vector) return int1530_t;
subtype uint1531_t is unsigned(1530 downto 0);
constant uint1531_t_SLV_LEN : integer := 1531;
function uint1531_t_to_slv(x : uint1531_t) return std_logic_vector;
function slv_to_uint1531_t(x : std_logic_vector) return uint1531_t;
subtype int1531_t is signed(1530 downto 0);
constant int1531_t_SLV_LEN : integer := 1531;
function int1531_t_to_slv(x : int1531_t) return std_logic_vector;
function slv_to_int1531_t(x : std_logic_vector) return int1531_t;
subtype uint1532_t is unsigned(1531 downto 0);
constant uint1532_t_SLV_LEN : integer := 1532;
function uint1532_t_to_slv(x : uint1532_t) return std_logic_vector;
function slv_to_uint1532_t(x : std_logic_vector) return uint1532_t;
subtype int1532_t is signed(1531 downto 0);
constant int1532_t_SLV_LEN : integer := 1532;
function int1532_t_to_slv(x : int1532_t) return std_logic_vector;
function slv_to_int1532_t(x : std_logic_vector) return int1532_t;
subtype uint1533_t is unsigned(1532 downto 0);
constant uint1533_t_SLV_LEN : integer := 1533;
function uint1533_t_to_slv(x : uint1533_t) return std_logic_vector;
function slv_to_uint1533_t(x : std_logic_vector) return uint1533_t;
subtype int1533_t is signed(1532 downto 0);
constant int1533_t_SLV_LEN : integer := 1533;
function int1533_t_to_slv(x : int1533_t) return std_logic_vector;
function slv_to_int1533_t(x : std_logic_vector) return int1533_t;
subtype uint1534_t is unsigned(1533 downto 0);
constant uint1534_t_SLV_LEN : integer := 1534;
function uint1534_t_to_slv(x : uint1534_t) return std_logic_vector;
function slv_to_uint1534_t(x : std_logic_vector) return uint1534_t;
subtype int1534_t is signed(1533 downto 0);
constant int1534_t_SLV_LEN : integer := 1534;
function int1534_t_to_slv(x : int1534_t) return std_logic_vector;
function slv_to_int1534_t(x : std_logic_vector) return int1534_t;
subtype uint1535_t is unsigned(1534 downto 0);
constant uint1535_t_SLV_LEN : integer := 1535;
function uint1535_t_to_slv(x : uint1535_t) return std_logic_vector;
function slv_to_uint1535_t(x : std_logic_vector) return uint1535_t;
subtype int1535_t is signed(1534 downto 0);
constant int1535_t_SLV_LEN : integer := 1535;
function int1535_t_to_slv(x : int1535_t) return std_logic_vector;
function slv_to_int1535_t(x : std_logic_vector) return int1535_t;
subtype uint1536_t is unsigned(1535 downto 0);
constant uint1536_t_SLV_LEN : integer := 1536;
function uint1536_t_to_slv(x : uint1536_t) return std_logic_vector;
function slv_to_uint1536_t(x : std_logic_vector) return uint1536_t;
subtype int1536_t is signed(1535 downto 0);
constant int1536_t_SLV_LEN : integer := 1536;
function int1536_t_to_slv(x : int1536_t) return std_logic_vector;
function slv_to_int1536_t(x : std_logic_vector) return int1536_t;
subtype uint1537_t is unsigned(1536 downto 0);
constant uint1537_t_SLV_LEN : integer := 1537;
function uint1537_t_to_slv(x : uint1537_t) return std_logic_vector;
function slv_to_uint1537_t(x : std_logic_vector) return uint1537_t;
subtype int1537_t is signed(1536 downto 0);
constant int1537_t_SLV_LEN : integer := 1537;
function int1537_t_to_slv(x : int1537_t) return std_logic_vector;
function slv_to_int1537_t(x : std_logic_vector) return int1537_t;
subtype uint1538_t is unsigned(1537 downto 0);
constant uint1538_t_SLV_LEN : integer := 1538;
function uint1538_t_to_slv(x : uint1538_t) return std_logic_vector;
function slv_to_uint1538_t(x : std_logic_vector) return uint1538_t;
subtype int1538_t is signed(1537 downto 0);
constant int1538_t_SLV_LEN : integer := 1538;
function int1538_t_to_slv(x : int1538_t) return std_logic_vector;
function slv_to_int1538_t(x : std_logic_vector) return int1538_t;
subtype uint1539_t is unsigned(1538 downto 0);
constant uint1539_t_SLV_LEN : integer := 1539;
function uint1539_t_to_slv(x : uint1539_t) return std_logic_vector;
function slv_to_uint1539_t(x : std_logic_vector) return uint1539_t;
subtype int1539_t is signed(1538 downto 0);
constant int1539_t_SLV_LEN : integer := 1539;
function int1539_t_to_slv(x : int1539_t) return std_logic_vector;
function slv_to_int1539_t(x : std_logic_vector) return int1539_t;
subtype uint1540_t is unsigned(1539 downto 0);
constant uint1540_t_SLV_LEN : integer := 1540;
function uint1540_t_to_slv(x : uint1540_t) return std_logic_vector;
function slv_to_uint1540_t(x : std_logic_vector) return uint1540_t;
subtype int1540_t is signed(1539 downto 0);
constant int1540_t_SLV_LEN : integer := 1540;
function int1540_t_to_slv(x : int1540_t) return std_logic_vector;
function slv_to_int1540_t(x : std_logic_vector) return int1540_t;
subtype uint1541_t is unsigned(1540 downto 0);
constant uint1541_t_SLV_LEN : integer := 1541;
function uint1541_t_to_slv(x : uint1541_t) return std_logic_vector;
function slv_to_uint1541_t(x : std_logic_vector) return uint1541_t;
subtype int1541_t is signed(1540 downto 0);
constant int1541_t_SLV_LEN : integer := 1541;
function int1541_t_to_slv(x : int1541_t) return std_logic_vector;
function slv_to_int1541_t(x : std_logic_vector) return int1541_t;
subtype uint1542_t is unsigned(1541 downto 0);
constant uint1542_t_SLV_LEN : integer := 1542;
function uint1542_t_to_slv(x : uint1542_t) return std_logic_vector;
function slv_to_uint1542_t(x : std_logic_vector) return uint1542_t;
subtype int1542_t is signed(1541 downto 0);
constant int1542_t_SLV_LEN : integer := 1542;
function int1542_t_to_slv(x : int1542_t) return std_logic_vector;
function slv_to_int1542_t(x : std_logic_vector) return int1542_t;
subtype uint1543_t is unsigned(1542 downto 0);
constant uint1543_t_SLV_LEN : integer := 1543;
function uint1543_t_to_slv(x : uint1543_t) return std_logic_vector;
function slv_to_uint1543_t(x : std_logic_vector) return uint1543_t;
subtype int1543_t is signed(1542 downto 0);
constant int1543_t_SLV_LEN : integer := 1543;
function int1543_t_to_slv(x : int1543_t) return std_logic_vector;
function slv_to_int1543_t(x : std_logic_vector) return int1543_t;
subtype uint1544_t is unsigned(1543 downto 0);
constant uint1544_t_SLV_LEN : integer := 1544;
function uint1544_t_to_slv(x : uint1544_t) return std_logic_vector;
function slv_to_uint1544_t(x : std_logic_vector) return uint1544_t;
subtype int1544_t is signed(1543 downto 0);
constant int1544_t_SLV_LEN : integer := 1544;
function int1544_t_to_slv(x : int1544_t) return std_logic_vector;
function slv_to_int1544_t(x : std_logic_vector) return int1544_t;
subtype uint1545_t is unsigned(1544 downto 0);
constant uint1545_t_SLV_LEN : integer := 1545;
function uint1545_t_to_slv(x : uint1545_t) return std_logic_vector;
function slv_to_uint1545_t(x : std_logic_vector) return uint1545_t;
subtype int1545_t is signed(1544 downto 0);
constant int1545_t_SLV_LEN : integer := 1545;
function int1545_t_to_slv(x : int1545_t) return std_logic_vector;
function slv_to_int1545_t(x : std_logic_vector) return int1545_t;
subtype uint1546_t is unsigned(1545 downto 0);
constant uint1546_t_SLV_LEN : integer := 1546;
function uint1546_t_to_slv(x : uint1546_t) return std_logic_vector;
function slv_to_uint1546_t(x : std_logic_vector) return uint1546_t;
subtype int1546_t is signed(1545 downto 0);
constant int1546_t_SLV_LEN : integer := 1546;
function int1546_t_to_slv(x : int1546_t) return std_logic_vector;
function slv_to_int1546_t(x : std_logic_vector) return int1546_t;
subtype uint1547_t is unsigned(1546 downto 0);
constant uint1547_t_SLV_LEN : integer := 1547;
function uint1547_t_to_slv(x : uint1547_t) return std_logic_vector;
function slv_to_uint1547_t(x : std_logic_vector) return uint1547_t;
subtype int1547_t is signed(1546 downto 0);
constant int1547_t_SLV_LEN : integer := 1547;
function int1547_t_to_slv(x : int1547_t) return std_logic_vector;
function slv_to_int1547_t(x : std_logic_vector) return int1547_t;
subtype uint1548_t is unsigned(1547 downto 0);
constant uint1548_t_SLV_LEN : integer := 1548;
function uint1548_t_to_slv(x : uint1548_t) return std_logic_vector;
function slv_to_uint1548_t(x : std_logic_vector) return uint1548_t;
subtype int1548_t is signed(1547 downto 0);
constant int1548_t_SLV_LEN : integer := 1548;
function int1548_t_to_slv(x : int1548_t) return std_logic_vector;
function slv_to_int1548_t(x : std_logic_vector) return int1548_t;
subtype uint1549_t is unsigned(1548 downto 0);
constant uint1549_t_SLV_LEN : integer := 1549;
function uint1549_t_to_slv(x : uint1549_t) return std_logic_vector;
function slv_to_uint1549_t(x : std_logic_vector) return uint1549_t;
subtype int1549_t is signed(1548 downto 0);
constant int1549_t_SLV_LEN : integer := 1549;
function int1549_t_to_slv(x : int1549_t) return std_logic_vector;
function slv_to_int1549_t(x : std_logic_vector) return int1549_t;
subtype uint1550_t is unsigned(1549 downto 0);
constant uint1550_t_SLV_LEN : integer := 1550;
function uint1550_t_to_slv(x : uint1550_t) return std_logic_vector;
function slv_to_uint1550_t(x : std_logic_vector) return uint1550_t;
subtype int1550_t is signed(1549 downto 0);
constant int1550_t_SLV_LEN : integer := 1550;
function int1550_t_to_slv(x : int1550_t) return std_logic_vector;
function slv_to_int1550_t(x : std_logic_vector) return int1550_t;
subtype uint1551_t is unsigned(1550 downto 0);
constant uint1551_t_SLV_LEN : integer := 1551;
function uint1551_t_to_slv(x : uint1551_t) return std_logic_vector;
function slv_to_uint1551_t(x : std_logic_vector) return uint1551_t;
subtype int1551_t is signed(1550 downto 0);
constant int1551_t_SLV_LEN : integer := 1551;
function int1551_t_to_slv(x : int1551_t) return std_logic_vector;
function slv_to_int1551_t(x : std_logic_vector) return int1551_t;
subtype uint1552_t is unsigned(1551 downto 0);
constant uint1552_t_SLV_LEN : integer := 1552;
function uint1552_t_to_slv(x : uint1552_t) return std_logic_vector;
function slv_to_uint1552_t(x : std_logic_vector) return uint1552_t;
subtype int1552_t is signed(1551 downto 0);
constant int1552_t_SLV_LEN : integer := 1552;
function int1552_t_to_slv(x : int1552_t) return std_logic_vector;
function slv_to_int1552_t(x : std_logic_vector) return int1552_t;
subtype uint1553_t is unsigned(1552 downto 0);
constant uint1553_t_SLV_LEN : integer := 1553;
function uint1553_t_to_slv(x : uint1553_t) return std_logic_vector;
function slv_to_uint1553_t(x : std_logic_vector) return uint1553_t;
subtype int1553_t is signed(1552 downto 0);
constant int1553_t_SLV_LEN : integer := 1553;
function int1553_t_to_slv(x : int1553_t) return std_logic_vector;
function slv_to_int1553_t(x : std_logic_vector) return int1553_t;
subtype uint1554_t is unsigned(1553 downto 0);
constant uint1554_t_SLV_LEN : integer := 1554;
function uint1554_t_to_slv(x : uint1554_t) return std_logic_vector;
function slv_to_uint1554_t(x : std_logic_vector) return uint1554_t;
subtype int1554_t is signed(1553 downto 0);
constant int1554_t_SLV_LEN : integer := 1554;
function int1554_t_to_slv(x : int1554_t) return std_logic_vector;
function slv_to_int1554_t(x : std_logic_vector) return int1554_t;
subtype uint1555_t is unsigned(1554 downto 0);
constant uint1555_t_SLV_LEN : integer := 1555;
function uint1555_t_to_slv(x : uint1555_t) return std_logic_vector;
function slv_to_uint1555_t(x : std_logic_vector) return uint1555_t;
subtype int1555_t is signed(1554 downto 0);
constant int1555_t_SLV_LEN : integer := 1555;
function int1555_t_to_slv(x : int1555_t) return std_logic_vector;
function slv_to_int1555_t(x : std_logic_vector) return int1555_t;
subtype uint1556_t is unsigned(1555 downto 0);
constant uint1556_t_SLV_LEN : integer := 1556;
function uint1556_t_to_slv(x : uint1556_t) return std_logic_vector;
function slv_to_uint1556_t(x : std_logic_vector) return uint1556_t;
subtype int1556_t is signed(1555 downto 0);
constant int1556_t_SLV_LEN : integer := 1556;
function int1556_t_to_slv(x : int1556_t) return std_logic_vector;
function slv_to_int1556_t(x : std_logic_vector) return int1556_t;
subtype uint1557_t is unsigned(1556 downto 0);
constant uint1557_t_SLV_LEN : integer := 1557;
function uint1557_t_to_slv(x : uint1557_t) return std_logic_vector;
function slv_to_uint1557_t(x : std_logic_vector) return uint1557_t;
subtype int1557_t is signed(1556 downto 0);
constant int1557_t_SLV_LEN : integer := 1557;
function int1557_t_to_slv(x : int1557_t) return std_logic_vector;
function slv_to_int1557_t(x : std_logic_vector) return int1557_t;
subtype uint1558_t is unsigned(1557 downto 0);
constant uint1558_t_SLV_LEN : integer := 1558;
function uint1558_t_to_slv(x : uint1558_t) return std_logic_vector;
function slv_to_uint1558_t(x : std_logic_vector) return uint1558_t;
subtype int1558_t is signed(1557 downto 0);
constant int1558_t_SLV_LEN : integer := 1558;
function int1558_t_to_slv(x : int1558_t) return std_logic_vector;
function slv_to_int1558_t(x : std_logic_vector) return int1558_t;
subtype uint1559_t is unsigned(1558 downto 0);
constant uint1559_t_SLV_LEN : integer := 1559;
function uint1559_t_to_slv(x : uint1559_t) return std_logic_vector;
function slv_to_uint1559_t(x : std_logic_vector) return uint1559_t;
subtype int1559_t is signed(1558 downto 0);
constant int1559_t_SLV_LEN : integer := 1559;
function int1559_t_to_slv(x : int1559_t) return std_logic_vector;
function slv_to_int1559_t(x : std_logic_vector) return int1559_t;
subtype uint1560_t is unsigned(1559 downto 0);
constant uint1560_t_SLV_LEN : integer := 1560;
function uint1560_t_to_slv(x : uint1560_t) return std_logic_vector;
function slv_to_uint1560_t(x : std_logic_vector) return uint1560_t;
subtype int1560_t is signed(1559 downto 0);
constant int1560_t_SLV_LEN : integer := 1560;
function int1560_t_to_slv(x : int1560_t) return std_logic_vector;
function slv_to_int1560_t(x : std_logic_vector) return int1560_t;
subtype uint1561_t is unsigned(1560 downto 0);
constant uint1561_t_SLV_LEN : integer := 1561;
function uint1561_t_to_slv(x : uint1561_t) return std_logic_vector;
function slv_to_uint1561_t(x : std_logic_vector) return uint1561_t;
subtype int1561_t is signed(1560 downto 0);
constant int1561_t_SLV_LEN : integer := 1561;
function int1561_t_to_slv(x : int1561_t) return std_logic_vector;
function slv_to_int1561_t(x : std_logic_vector) return int1561_t;
subtype uint1562_t is unsigned(1561 downto 0);
constant uint1562_t_SLV_LEN : integer := 1562;
function uint1562_t_to_slv(x : uint1562_t) return std_logic_vector;
function slv_to_uint1562_t(x : std_logic_vector) return uint1562_t;
subtype int1562_t is signed(1561 downto 0);
constant int1562_t_SLV_LEN : integer := 1562;
function int1562_t_to_slv(x : int1562_t) return std_logic_vector;
function slv_to_int1562_t(x : std_logic_vector) return int1562_t;
subtype uint1563_t is unsigned(1562 downto 0);
constant uint1563_t_SLV_LEN : integer := 1563;
function uint1563_t_to_slv(x : uint1563_t) return std_logic_vector;
function slv_to_uint1563_t(x : std_logic_vector) return uint1563_t;
subtype int1563_t is signed(1562 downto 0);
constant int1563_t_SLV_LEN : integer := 1563;
function int1563_t_to_slv(x : int1563_t) return std_logic_vector;
function slv_to_int1563_t(x : std_logic_vector) return int1563_t;
subtype uint1564_t is unsigned(1563 downto 0);
constant uint1564_t_SLV_LEN : integer := 1564;
function uint1564_t_to_slv(x : uint1564_t) return std_logic_vector;
function slv_to_uint1564_t(x : std_logic_vector) return uint1564_t;
subtype int1564_t is signed(1563 downto 0);
constant int1564_t_SLV_LEN : integer := 1564;
function int1564_t_to_slv(x : int1564_t) return std_logic_vector;
function slv_to_int1564_t(x : std_logic_vector) return int1564_t;
subtype uint1565_t is unsigned(1564 downto 0);
constant uint1565_t_SLV_LEN : integer := 1565;
function uint1565_t_to_slv(x : uint1565_t) return std_logic_vector;
function slv_to_uint1565_t(x : std_logic_vector) return uint1565_t;
subtype int1565_t is signed(1564 downto 0);
constant int1565_t_SLV_LEN : integer := 1565;
function int1565_t_to_slv(x : int1565_t) return std_logic_vector;
function slv_to_int1565_t(x : std_logic_vector) return int1565_t;
subtype uint1566_t is unsigned(1565 downto 0);
constant uint1566_t_SLV_LEN : integer := 1566;
function uint1566_t_to_slv(x : uint1566_t) return std_logic_vector;
function slv_to_uint1566_t(x : std_logic_vector) return uint1566_t;
subtype int1566_t is signed(1565 downto 0);
constant int1566_t_SLV_LEN : integer := 1566;
function int1566_t_to_slv(x : int1566_t) return std_logic_vector;
function slv_to_int1566_t(x : std_logic_vector) return int1566_t;
subtype uint1567_t is unsigned(1566 downto 0);
constant uint1567_t_SLV_LEN : integer := 1567;
function uint1567_t_to_slv(x : uint1567_t) return std_logic_vector;
function slv_to_uint1567_t(x : std_logic_vector) return uint1567_t;
subtype int1567_t is signed(1566 downto 0);
constant int1567_t_SLV_LEN : integer := 1567;
function int1567_t_to_slv(x : int1567_t) return std_logic_vector;
function slv_to_int1567_t(x : std_logic_vector) return int1567_t;
subtype uint1568_t is unsigned(1567 downto 0);
constant uint1568_t_SLV_LEN : integer := 1568;
function uint1568_t_to_slv(x : uint1568_t) return std_logic_vector;
function slv_to_uint1568_t(x : std_logic_vector) return uint1568_t;
subtype int1568_t is signed(1567 downto 0);
constant int1568_t_SLV_LEN : integer := 1568;
function int1568_t_to_slv(x : int1568_t) return std_logic_vector;
function slv_to_int1568_t(x : std_logic_vector) return int1568_t;
subtype uint1569_t is unsigned(1568 downto 0);
constant uint1569_t_SLV_LEN : integer := 1569;
function uint1569_t_to_slv(x : uint1569_t) return std_logic_vector;
function slv_to_uint1569_t(x : std_logic_vector) return uint1569_t;
subtype int1569_t is signed(1568 downto 0);
constant int1569_t_SLV_LEN : integer := 1569;
function int1569_t_to_slv(x : int1569_t) return std_logic_vector;
function slv_to_int1569_t(x : std_logic_vector) return int1569_t;
subtype uint1570_t is unsigned(1569 downto 0);
constant uint1570_t_SLV_LEN : integer := 1570;
function uint1570_t_to_slv(x : uint1570_t) return std_logic_vector;
function slv_to_uint1570_t(x : std_logic_vector) return uint1570_t;
subtype int1570_t is signed(1569 downto 0);
constant int1570_t_SLV_LEN : integer := 1570;
function int1570_t_to_slv(x : int1570_t) return std_logic_vector;
function slv_to_int1570_t(x : std_logic_vector) return int1570_t;
subtype uint1571_t is unsigned(1570 downto 0);
constant uint1571_t_SLV_LEN : integer := 1571;
function uint1571_t_to_slv(x : uint1571_t) return std_logic_vector;
function slv_to_uint1571_t(x : std_logic_vector) return uint1571_t;
subtype int1571_t is signed(1570 downto 0);
constant int1571_t_SLV_LEN : integer := 1571;
function int1571_t_to_slv(x : int1571_t) return std_logic_vector;
function slv_to_int1571_t(x : std_logic_vector) return int1571_t;
subtype uint1572_t is unsigned(1571 downto 0);
constant uint1572_t_SLV_LEN : integer := 1572;
function uint1572_t_to_slv(x : uint1572_t) return std_logic_vector;
function slv_to_uint1572_t(x : std_logic_vector) return uint1572_t;
subtype int1572_t is signed(1571 downto 0);
constant int1572_t_SLV_LEN : integer := 1572;
function int1572_t_to_slv(x : int1572_t) return std_logic_vector;
function slv_to_int1572_t(x : std_logic_vector) return int1572_t;
subtype uint1573_t is unsigned(1572 downto 0);
constant uint1573_t_SLV_LEN : integer := 1573;
function uint1573_t_to_slv(x : uint1573_t) return std_logic_vector;
function slv_to_uint1573_t(x : std_logic_vector) return uint1573_t;
subtype int1573_t is signed(1572 downto 0);
constant int1573_t_SLV_LEN : integer := 1573;
function int1573_t_to_slv(x : int1573_t) return std_logic_vector;
function slv_to_int1573_t(x : std_logic_vector) return int1573_t;
subtype uint1574_t is unsigned(1573 downto 0);
constant uint1574_t_SLV_LEN : integer := 1574;
function uint1574_t_to_slv(x : uint1574_t) return std_logic_vector;
function slv_to_uint1574_t(x : std_logic_vector) return uint1574_t;
subtype int1574_t is signed(1573 downto 0);
constant int1574_t_SLV_LEN : integer := 1574;
function int1574_t_to_slv(x : int1574_t) return std_logic_vector;
function slv_to_int1574_t(x : std_logic_vector) return int1574_t;
subtype uint1575_t is unsigned(1574 downto 0);
constant uint1575_t_SLV_LEN : integer := 1575;
function uint1575_t_to_slv(x : uint1575_t) return std_logic_vector;
function slv_to_uint1575_t(x : std_logic_vector) return uint1575_t;
subtype int1575_t is signed(1574 downto 0);
constant int1575_t_SLV_LEN : integer := 1575;
function int1575_t_to_slv(x : int1575_t) return std_logic_vector;
function slv_to_int1575_t(x : std_logic_vector) return int1575_t;
subtype uint1576_t is unsigned(1575 downto 0);
constant uint1576_t_SLV_LEN : integer := 1576;
function uint1576_t_to_slv(x : uint1576_t) return std_logic_vector;
function slv_to_uint1576_t(x : std_logic_vector) return uint1576_t;
subtype int1576_t is signed(1575 downto 0);
constant int1576_t_SLV_LEN : integer := 1576;
function int1576_t_to_slv(x : int1576_t) return std_logic_vector;
function slv_to_int1576_t(x : std_logic_vector) return int1576_t;
subtype uint1577_t is unsigned(1576 downto 0);
constant uint1577_t_SLV_LEN : integer := 1577;
function uint1577_t_to_slv(x : uint1577_t) return std_logic_vector;
function slv_to_uint1577_t(x : std_logic_vector) return uint1577_t;
subtype int1577_t is signed(1576 downto 0);
constant int1577_t_SLV_LEN : integer := 1577;
function int1577_t_to_slv(x : int1577_t) return std_logic_vector;
function slv_to_int1577_t(x : std_logic_vector) return int1577_t;
subtype uint1578_t is unsigned(1577 downto 0);
constant uint1578_t_SLV_LEN : integer := 1578;
function uint1578_t_to_slv(x : uint1578_t) return std_logic_vector;
function slv_to_uint1578_t(x : std_logic_vector) return uint1578_t;
subtype int1578_t is signed(1577 downto 0);
constant int1578_t_SLV_LEN : integer := 1578;
function int1578_t_to_slv(x : int1578_t) return std_logic_vector;
function slv_to_int1578_t(x : std_logic_vector) return int1578_t;
subtype uint1579_t is unsigned(1578 downto 0);
constant uint1579_t_SLV_LEN : integer := 1579;
function uint1579_t_to_slv(x : uint1579_t) return std_logic_vector;
function slv_to_uint1579_t(x : std_logic_vector) return uint1579_t;
subtype int1579_t is signed(1578 downto 0);
constant int1579_t_SLV_LEN : integer := 1579;
function int1579_t_to_slv(x : int1579_t) return std_logic_vector;
function slv_to_int1579_t(x : std_logic_vector) return int1579_t;
subtype uint1580_t is unsigned(1579 downto 0);
constant uint1580_t_SLV_LEN : integer := 1580;
function uint1580_t_to_slv(x : uint1580_t) return std_logic_vector;
function slv_to_uint1580_t(x : std_logic_vector) return uint1580_t;
subtype int1580_t is signed(1579 downto 0);
constant int1580_t_SLV_LEN : integer := 1580;
function int1580_t_to_slv(x : int1580_t) return std_logic_vector;
function slv_to_int1580_t(x : std_logic_vector) return int1580_t;
subtype uint1581_t is unsigned(1580 downto 0);
constant uint1581_t_SLV_LEN : integer := 1581;
function uint1581_t_to_slv(x : uint1581_t) return std_logic_vector;
function slv_to_uint1581_t(x : std_logic_vector) return uint1581_t;
subtype int1581_t is signed(1580 downto 0);
constant int1581_t_SLV_LEN : integer := 1581;
function int1581_t_to_slv(x : int1581_t) return std_logic_vector;
function slv_to_int1581_t(x : std_logic_vector) return int1581_t;
subtype uint1582_t is unsigned(1581 downto 0);
constant uint1582_t_SLV_LEN : integer := 1582;
function uint1582_t_to_slv(x : uint1582_t) return std_logic_vector;
function slv_to_uint1582_t(x : std_logic_vector) return uint1582_t;
subtype int1582_t is signed(1581 downto 0);
constant int1582_t_SLV_LEN : integer := 1582;
function int1582_t_to_slv(x : int1582_t) return std_logic_vector;
function slv_to_int1582_t(x : std_logic_vector) return int1582_t;
subtype uint1583_t is unsigned(1582 downto 0);
constant uint1583_t_SLV_LEN : integer := 1583;
function uint1583_t_to_slv(x : uint1583_t) return std_logic_vector;
function slv_to_uint1583_t(x : std_logic_vector) return uint1583_t;
subtype int1583_t is signed(1582 downto 0);
constant int1583_t_SLV_LEN : integer := 1583;
function int1583_t_to_slv(x : int1583_t) return std_logic_vector;
function slv_to_int1583_t(x : std_logic_vector) return int1583_t;
subtype uint1584_t is unsigned(1583 downto 0);
constant uint1584_t_SLV_LEN : integer := 1584;
function uint1584_t_to_slv(x : uint1584_t) return std_logic_vector;
function slv_to_uint1584_t(x : std_logic_vector) return uint1584_t;
subtype int1584_t is signed(1583 downto 0);
constant int1584_t_SLV_LEN : integer := 1584;
function int1584_t_to_slv(x : int1584_t) return std_logic_vector;
function slv_to_int1584_t(x : std_logic_vector) return int1584_t;
subtype uint1585_t is unsigned(1584 downto 0);
constant uint1585_t_SLV_LEN : integer := 1585;
function uint1585_t_to_slv(x : uint1585_t) return std_logic_vector;
function slv_to_uint1585_t(x : std_logic_vector) return uint1585_t;
subtype int1585_t is signed(1584 downto 0);
constant int1585_t_SLV_LEN : integer := 1585;
function int1585_t_to_slv(x : int1585_t) return std_logic_vector;
function slv_to_int1585_t(x : std_logic_vector) return int1585_t;
subtype uint1586_t is unsigned(1585 downto 0);
constant uint1586_t_SLV_LEN : integer := 1586;
function uint1586_t_to_slv(x : uint1586_t) return std_logic_vector;
function slv_to_uint1586_t(x : std_logic_vector) return uint1586_t;
subtype int1586_t is signed(1585 downto 0);
constant int1586_t_SLV_LEN : integer := 1586;
function int1586_t_to_slv(x : int1586_t) return std_logic_vector;
function slv_to_int1586_t(x : std_logic_vector) return int1586_t;
subtype uint1587_t is unsigned(1586 downto 0);
constant uint1587_t_SLV_LEN : integer := 1587;
function uint1587_t_to_slv(x : uint1587_t) return std_logic_vector;
function slv_to_uint1587_t(x : std_logic_vector) return uint1587_t;
subtype int1587_t is signed(1586 downto 0);
constant int1587_t_SLV_LEN : integer := 1587;
function int1587_t_to_slv(x : int1587_t) return std_logic_vector;
function slv_to_int1587_t(x : std_logic_vector) return int1587_t;
subtype uint1588_t is unsigned(1587 downto 0);
constant uint1588_t_SLV_LEN : integer := 1588;
function uint1588_t_to_slv(x : uint1588_t) return std_logic_vector;
function slv_to_uint1588_t(x : std_logic_vector) return uint1588_t;
subtype int1588_t is signed(1587 downto 0);
constant int1588_t_SLV_LEN : integer := 1588;
function int1588_t_to_slv(x : int1588_t) return std_logic_vector;
function slv_to_int1588_t(x : std_logic_vector) return int1588_t;
subtype uint1589_t is unsigned(1588 downto 0);
constant uint1589_t_SLV_LEN : integer := 1589;
function uint1589_t_to_slv(x : uint1589_t) return std_logic_vector;
function slv_to_uint1589_t(x : std_logic_vector) return uint1589_t;
subtype int1589_t is signed(1588 downto 0);
constant int1589_t_SLV_LEN : integer := 1589;
function int1589_t_to_slv(x : int1589_t) return std_logic_vector;
function slv_to_int1589_t(x : std_logic_vector) return int1589_t;
subtype uint1590_t is unsigned(1589 downto 0);
constant uint1590_t_SLV_LEN : integer := 1590;
function uint1590_t_to_slv(x : uint1590_t) return std_logic_vector;
function slv_to_uint1590_t(x : std_logic_vector) return uint1590_t;
subtype int1590_t is signed(1589 downto 0);
constant int1590_t_SLV_LEN : integer := 1590;
function int1590_t_to_slv(x : int1590_t) return std_logic_vector;
function slv_to_int1590_t(x : std_logic_vector) return int1590_t;
subtype uint1591_t is unsigned(1590 downto 0);
constant uint1591_t_SLV_LEN : integer := 1591;
function uint1591_t_to_slv(x : uint1591_t) return std_logic_vector;
function slv_to_uint1591_t(x : std_logic_vector) return uint1591_t;
subtype int1591_t is signed(1590 downto 0);
constant int1591_t_SLV_LEN : integer := 1591;
function int1591_t_to_slv(x : int1591_t) return std_logic_vector;
function slv_to_int1591_t(x : std_logic_vector) return int1591_t;
subtype uint1592_t is unsigned(1591 downto 0);
constant uint1592_t_SLV_LEN : integer := 1592;
function uint1592_t_to_slv(x : uint1592_t) return std_logic_vector;
function slv_to_uint1592_t(x : std_logic_vector) return uint1592_t;
subtype int1592_t is signed(1591 downto 0);
constant int1592_t_SLV_LEN : integer := 1592;
function int1592_t_to_slv(x : int1592_t) return std_logic_vector;
function slv_to_int1592_t(x : std_logic_vector) return int1592_t;
subtype uint1593_t is unsigned(1592 downto 0);
constant uint1593_t_SLV_LEN : integer := 1593;
function uint1593_t_to_slv(x : uint1593_t) return std_logic_vector;
function slv_to_uint1593_t(x : std_logic_vector) return uint1593_t;
subtype int1593_t is signed(1592 downto 0);
constant int1593_t_SLV_LEN : integer := 1593;
function int1593_t_to_slv(x : int1593_t) return std_logic_vector;
function slv_to_int1593_t(x : std_logic_vector) return int1593_t;
subtype uint1594_t is unsigned(1593 downto 0);
constant uint1594_t_SLV_LEN : integer := 1594;
function uint1594_t_to_slv(x : uint1594_t) return std_logic_vector;
function slv_to_uint1594_t(x : std_logic_vector) return uint1594_t;
subtype int1594_t is signed(1593 downto 0);
constant int1594_t_SLV_LEN : integer := 1594;
function int1594_t_to_slv(x : int1594_t) return std_logic_vector;
function slv_to_int1594_t(x : std_logic_vector) return int1594_t;
subtype uint1595_t is unsigned(1594 downto 0);
constant uint1595_t_SLV_LEN : integer := 1595;
function uint1595_t_to_slv(x : uint1595_t) return std_logic_vector;
function slv_to_uint1595_t(x : std_logic_vector) return uint1595_t;
subtype int1595_t is signed(1594 downto 0);
constant int1595_t_SLV_LEN : integer := 1595;
function int1595_t_to_slv(x : int1595_t) return std_logic_vector;
function slv_to_int1595_t(x : std_logic_vector) return int1595_t;
subtype uint1596_t is unsigned(1595 downto 0);
constant uint1596_t_SLV_LEN : integer := 1596;
function uint1596_t_to_slv(x : uint1596_t) return std_logic_vector;
function slv_to_uint1596_t(x : std_logic_vector) return uint1596_t;
subtype int1596_t is signed(1595 downto 0);
constant int1596_t_SLV_LEN : integer := 1596;
function int1596_t_to_slv(x : int1596_t) return std_logic_vector;
function slv_to_int1596_t(x : std_logic_vector) return int1596_t;
subtype uint1597_t is unsigned(1596 downto 0);
constant uint1597_t_SLV_LEN : integer := 1597;
function uint1597_t_to_slv(x : uint1597_t) return std_logic_vector;
function slv_to_uint1597_t(x : std_logic_vector) return uint1597_t;
subtype int1597_t is signed(1596 downto 0);
constant int1597_t_SLV_LEN : integer := 1597;
function int1597_t_to_slv(x : int1597_t) return std_logic_vector;
function slv_to_int1597_t(x : std_logic_vector) return int1597_t;
subtype uint1598_t is unsigned(1597 downto 0);
constant uint1598_t_SLV_LEN : integer := 1598;
function uint1598_t_to_slv(x : uint1598_t) return std_logic_vector;
function slv_to_uint1598_t(x : std_logic_vector) return uint1598_t;
subtype int1598_t is signed(1597 downto 0);
constant int1598_t_SLV_LEN : integer := 1598;
function int1598_t_to_slv(x : int1598_t) return std_logic_vector;
function slv_to_int1598_t(x : std_logic_vector) return int1598_t;
subtype uint1599_t is unsigned(1598 downto 0);
constant uint1599_t_SLV_LEN : integer := 1599;
function uint1599_t_to_slv(x : uint1599_t) return std_logic_vector;
function slv_to_uint1599_t(x : std_logic_vector) return uint1599_t;
subtype int1599_t is signed(1598 downto 0);
constant int1599_t_SLV_LEN : integer := 1599;
function int1599_t_to_slv(x : int1599_t) return std_logic_vector;
function slv_to_int1599_t(x : std_logic_vector) return int1599_t;
subtype uint1600_t is unsigned(1599 downto 0);
constant uint1600_t_SLV_LEN : integer := 1600;
function uint1600_t_to_slv(x : uint1600_t) return std_logic_vector;
function slv_to_uint1600_t(x : std_logic_vector) return uint1600_t;
subtype int1600_t is signed(1599 downto 0);
constant int1600_t_SLV_LEN : integer := 1600;
function int1600_t_to_slv(x : int1600_t) return std_logic_vector;
function slv_to_int1600_t(x : std_logic_vector) return int1600_t;
subtype uint1601_t is unsigned(1600 downto 0);
constant uint1601_t_SLV_LEN : integer := 1601;
function uint1601_t_to_slv(x : uint1601_t) return std_logic_vector;
function slv_to_uint1601_t(x : std_logic_vector) return uint1601_t;
subtype int1601_t is signed(1600 downto 0);
constant int1601_t_SLV_LEN : integer := 1601;
function int1601_t_to_slv(x : int1601_t) return std_logic_vector;
function slv_to_int1601_t(x : std_logic_vector) return int1601_t;
subtype uint1602_t is unsigned(1601 downto 0);
constant uint1602_t_SLV_LEN : integer := 1602;
function uint1602_t_to_slv(x : uint1602_t) return std_logic_vector;
function slv_to_uint1602_t(x : std_logic_vector) return uint1602_t;
subtype int1602_t is signed(1601 downto 0);
constant int1602_t_SLV_LEN : integer := 1602;
function int1602_t_to_slv(x : int1602_t) return std_logic_vector;
function slv_to_int1602_t(x : std_logic_vector) return int1602_t;
subtype uint1603_t is unsigned(1602 downto 0);
constant uint1603_t_SLV_LEN : integer := 1603;
function uint1603_t_to_slv(x : uint1603_t) return std_logic_vector;
function slv_to_uint1603_t(x : std_logic_vector) return uint1603_t;
subtype int1603_t is signed(1602 downto 0);
constant int1603_t_SLV_LEN : integer := 1603;
function int1603_t_to_slv(x : int1603_t) return std_logic_vector;
function slv_to_int1603_t(x : std_logic_vector) return int1603_t;
subtype uint1604_t is unsigned(1603 downto 0);
constant uint1604_t_SLV_LEN : integer := 1604;
function uint1604_t_to_slv(x : uint1604_t) return std_logic_vector;
function slv_to_uint1604_t(x : std_logic_vector) return uint1604_t;
subtype int1604_t is signed(1603 downto 0);
constant int1604_t_SLV_LEN : integer := 1604;
function int1604_t_to_slv(x : int1604_t) return std_logic_vector;
function slv_to_int1604_t(x : std_logic_vector) return int1604_t;
subtype uint1605_t is unsigned(1604 downto 0);
constant uint1605_t_SLV_LEN : integer := 1605;
function uint1605_t_to_slv(x : uint1605_t) return std_logic_vector;
function slv_to_uint1605_t(x : std_logic_vector) return uint1605_t;
subtype int1605_t is signed(1604 downto 0);
constant int1605_t_SLV_LEN : integer := 1605;
function int1605_t_to_slv(x : int1605_t) return std_logic_vector;
function slv_to_int1605_t(x : std_logic_vector) return int1605_t;
subtype uint1606_t is unsigned(1605 downto 0);
constant uint1606_t_SLV_LEN : integer := 1606;
function uint1606_t_to_slv(x : uint1606_t) return std_logic_vector;
function slv_to_uint1606_t(x : std_logic_vector) return uint1606_t;
subtype int1606_t is signed(1605 downto 0);
constant int1606_t_SLV_LEN : integer := 1606;
function int1606_t_to_slv(x : int1606_t) return std_logic_vector;
function slv_to_int1606_t(x : std_logic_vector) return int1606_t;
subtype uint1607_t is unsigned(1606 downto 0);
constant uint1607_t_SLV_LEN : integer := 1607;
function uint1607_t_to_slv(x : uint1607_t) return std_logic_vector;
function slv_to_uint1607_t(x : std_logic_vector) return uint1607_t;
subtype int1607_t is signed(1606 downto 0);
constant int1607_t_SLV_LEN : integer := 1607;
function int1607_t_to_slv(x : int1607_t) return std_logic_vector;
function slv_to_int1607_t(x : std_logic_vector) return int1607_t;
subtype uint1608_t is unsigned(1607 downto 0);
constant uint1608_t_SLV_LEN : integer := 1608;
function uint1608_t_to_slv(x : uint1608_t) return std_logic_vector;
function slv_to_uint1608_t(x : std_logic_vector) return uint1608_t;
subtype int1608_t is signed(1607 downto 0);
constant int1608_t_SLV_LEN : integer := 1608;
function int1608_t_to_slv(x : int1608_t) return std_logic_vector;
function slv_to_int1608_t(x : std_logic_vector) return int1608_t;
subtype uint1609_t is unsigned(1608 downto 0);
constant uint1609_t_SLV_LEN : integer := 1609;
function uint1609_t_to_slv(x : uint1609_t) return std_logic_vector;
function slv_to_uint1609_t(x : std_logic_vector) return uint1609_t;
subtype int1609_t is signed(1608 downto 0);
constant int1609_t_SLV_LEN : integer := 1609;
function int1609_t_to_slv(x : int1609_t) return std_logic_vector;
function slv_to_int1609_t(x : std_logic_vector) return int1609_t;
subtype uint1610_t is unsigned(1609 downto 0);
constant uint1610_t_SLV_LEN : integer := 1610;
function uint1610_t_to_slv(x : uint1610_t) return std_logic_vector;
function slv_to_uint1610_t(x : std_logic_vector) return uint1610_t;
subtype int1610_t is signed(1609 downto 0);
constant int1610_t_SLV_LEN : integer := 1610;
function int1610_t_to_slv(x : int1610_t) return std_logic_vector;
function slv_to_int1610_t(x : std_logic_vector) return int1610_t;
subtype uint1611_t is unsigned(1610 downto 0);
constant uint1611_t_SLV_LEN : integer := 1611;
function uint1611_t_to_slv(x : uint1611_t) return std_logic_vector;
function slv_to_uint1611_t(x : std_logic_vector) return uint1611_t;
subtype int1611_t is signed(1610 downto 0);
constant int1611_t_SLV_LEN : integer := 1611;
function int1611_t_to_slv(x : int1611_t) return std_logic_vector;
function slv_to_int1611_t(x : std_logic_vector) return int1611_t;
subtype uint1612_t is unsigned(1611 downto 0);
constant uint1612_t_SLV_LEN : integer := 1612;
function uint1612_t_to_slv(x : uint1612_t) return std_logic_vector;
function slv_to_uint1612_t(x : std_logic_vector) return uint1612_t;
subtype int1612_t is signed(1611 downto 0);
constant int1612_t_SLV_LEN : integer := 1612;
function int1612_t_to_slv(x : int1612_t) return std_logic_vector;
function slv_to_int1612_t(x : std_logic_vector) return int1612_t;
subtype uint1613_t is unsigned(1612 downto 0);
constant uint1613_t_SLV_LEN : integer := 1613;
function uint1613_t_to_slv(x : uint1613_t) return std_logic_vector;
function slv_to_uint1613_t(x : std_logic_vector) return uint1613_t;
subtype int1613_t is signed(1612 downto 0);
constant int1613_t_SLV_LEN : integer := 1613;
function int1613_t_to_slv(x : int1613_t) return std_logic_vector;
function slv_to_int1613_t(x : std_logic_vector) return int1613_t;
subtype uint1614_t is unsigned(1613 downto 0);
constant uint1614_t_SLV_LEN : integer := 1614;
function uint1614_t_to_slv(x : uint1614_t) return std_logic_vector;
function slv_to_uint1614_t(x : std_logic_vector) return uint1614_t;
subtype int1614_t is signed(1613 downto 0);
constant int1614_t_SLV_LEN : integer := 1614;
function int1614_t_to_slv(x : int1614_t) return std_logic_vector;
function slv_to_int1614_t(x : std_logic_vector) return int1614_t;
subtype uint1615_t is unsigned(1614 downto 0);
constant uint1615_t_SLV_LEN : integer := 1615;
function uint1615_t_to_slv(x : uint1615_t) return std_logic_vector;
function slv_to_uint1615_t(x : std_logic_vector) return uint1615_t;
subtype int1615_t is signed(1614 downto 0);
constant int1615_t_SLV_LEN : integer := 1615;
function int1615_t_to_slv(x : int1615_t) return std_logic_vector;
function slv_to_int1615_t(x : std_logic_vector) return int1615_t;
subtype uint1616_t is unsigned(1615 downto 0);
constant uint1616_t_SLV_LEN : integer := 1616;
function uint1616_t_to_slv(x : uint1616_t) return std_logic_vector;
function slv_to_uint1616_t(x : std_logic_vector) return uint1616_t;
subtype int1616_t is signed(1615 downto 0);
constant int1616_t_SLV_LEN : integer := 1616;
function int1616_t_to_slv(x : int1616_t) return std_logic_vector;
function slv_to_int1616_t(x : std_logic_vector) return int1616_t;
subtype uint1617_t is unsigned(1616 downto 0);
constant uint1617_t_SLV_LEN : integer := 1617;
function uint1617_t_to_slv(x : uint1617_t) return std_logic_vector;
function slv_to_uint1617_t(x : std_logic_vector) return uint1617_t;
subtype int1617_t is signed(1616 downto 0);
constant int1617_t_SLV_LEN : integer := 1617;
function int1617_t_to_slv(x : int1617_t) return std_logic_vector;
function slv_to_int1617_t(x : std_logic_vector) return int1617_t;
subtype uint1618_t is unsigned(1617 downto 0);
constant uint1618_t_SLV_LEN : integer := 1618;
function uint1618_t_to_slv(x : uint1618_t) return std_logic_vector;
function slv_to_uint1618_t(x : std_logic_vector) return uint1618_t;
subtype int1618_t is signed(1617 downto 0);
constant int1618_t_SLV_LEN : integer := 1618;
function int1618_t_to_slv(x : int1618_t) return std_logic_vector;
function slv_to_int1618_t(x : std_logic_vector) return int1618_t;
subtype uint1619_t is unsigned(1618 downto 0);
constant uint1619_t_SLV_LEN : integer := 1619;
function uint1619_t_to_slv(x : uint1619_t) return std_logic_vector;
function slv_to_uint1619_t(x : std_logic_vector) return uint1619_t;
subtype int1619_t is signed(1618 downto 0);
constant int1619_t_SLV_LEN : integer := 1619;
function int1619_t_to_slv(x : int1619_t) return std_logic_vector;
function slv_to_int1619_t(x : std_logic_vector) return int1619_t;
subtype uint1620_t is unsigned(1619 downto 0);
constant uint1620_t_SLV_LEN : integer := 1620;
function uint1620_t_to_slv(x : uint1620_t) return std_logic_vector;
function slv_to_uint1620_t(x : std_logic_vector) return uint1620_t;
subtype int1620_t is signed(1619 downto 0);
constant int1620_t_SLV_LEN : integer := 1620;
function int1620_t_to_slv(x : int1620_t) return std_logic_vector;
function slv_to_int1620_t(x : std_logic_vector) return int1620_t;
subtype uint1621_t is unsigned(1620 downto 0);
constant uint1621_t_SLV_LEN : integer := 1621;
function uint1621_t_to_slv(x : uint1621_t) return std_logic_vector;
function slv_to_uint1621_t(x : std_logic_vector) return uint1621_t;
subtype int1621_t is signed(1620 downto 0);
constant int1621_t_SLV_LEN : integer := 1621;
function int1621_t_to_slv(x : int1621_t) return std_logic_vector;
function slv_to_int1621_t(x : std_logic_vector) return int1621_t;
subtype uint1622_t is unsigned(1621 downto 0);
constant uint1622_t_SLV_LEN : integer := 1622;
function uint1622_t_to_slv(x : uint1622_t) return std_logic_vector;
function slv_to_uint1622_t(x : std_logic_vector) return uint1622_t;
subtype int1622_t is signed(1621 downto 0);
constant int1622_t_SLV_LEN : integer := 1622;
function int1622_t_to_slv(x : int1622_t) return std_logic_vector;
function slv_to_int1622_t(x : std_logic_vector) return int1622_t;
subtype uint1623_t is unsigned(1622 downto 0);
constant uint1623_t_SLV_LEN : integer := 1623;
function uint1623_t_to_slv(x : uint1623_t) return std_logic_vector;
function slv_to_uint1623_t(x : std_logic_vector) return uint1623_t;
subtype int1623_t is signed(1622 downto 0);
constant int1623_t_SLV_LEN : integer := 1623;
function int1623_t_to_slv(x : int1623_t) return std_logic_vector;
function slv_to_int1623_t(x : std_logic_vector) return int1623_t;
subtype uint1624_t is unsigned(1623 downto 0);
constant uint1624_t_SLV_LEN : integer := 1624;
function uint1624_t_to_slv(x : uint1624_t) return std_logic_vector;
function slv_to_uint1624_t(x : std_logic_vector) return uint1624_t;
subtype int1624_t is signed(1623 downto 0);
constant int1624_t_SLV_LEN : integer := 1624;
function int1624_t_to_slv(x : int1624_t) return std_logic_vector;
function slv_to_int1624_t(x : std_logic_vector) return int1624_t;
subtype uint1625_t is unsigned(1624 downto 0);
constant uint1625_t_SLV_LEN : integer := 1625;
function uint1625_t_to_slv(x : uint1625_t) return std_logic_vector;
function slv_to_uint1625_t(x : std_logic_vector) return uint1625_t;
subtype int1625_t is signed(1624 downto 0);
constant int1625_t_SLV_LEN : integer := 1625;
function int1625_t_to_slv(x : int1625_t) return std_logic_vector;
function slv_to_int1625_t(x : std_logic_vector) return int1625_t;
subtype uint1626_t is unsigned(1625 downto 0);
constant uint1626_t_SLV_LEN : integer := 1626;
function uint1626_t_to_slv(x : uint1626_t) return std_logic_vector;
function slv_to_uint1626_t(x : std_logic_vector) return uint1626_t;
subtype int1626_t is signed(1625 downto 0);
constant int1626_t_SLV_LEN : integer := 1626;
function int1626_t_to_slv(x : int1626_t) return std_logic_vector;
function slv_to_int1626_t(x : std_logic_vector) return int1626_t;
subtype uint1627_t is unsigned(1626 downto 0);
constant uint1627_t_SLV_LEN : integer := 1627;
function uint1627_t_to_slv(x : uint1627_t) return std_logic_vector;
function slv_to_uint1627_t(x : std_logic_vector) return uint1627_t;
subtype int1627_t is signed(1626 downto 0);
constant int1627_t_SLV_LEN : integer := 1627;
function int1627_t_to_slv(x : int1627_t) return std_logic_vector;
function slv_to_int1627_t(x : std_logic_vector) return int1627_t;
subtype uint1628_t is unsigned(1627 downto 0);
constant uint1628_t_SLV_LEN : integer := 1628;
function uint1628_t_to_slv(x : uint1628_t) return std_logic_vector;
function slv_to_uint1628_t(x : std_logic_vector) return uint1628_t;
subtype int1628_t is signed(1627 downto 0);
constant int1628_t_SLV_LEN : integer := 1628;
function int1628_t_to_slv(x : int1628_t) return std_logic_vector;
function slv_to_int1628_t(x : std_logic_vector) return int1628_t;
subtype uint1629_t is unsigned(1628 downto 0);
constant uint1629_t_SLV_LEN : integer := 1629;
function uint1629_t_to_slv(x : uint1629_t) return std_logic_vector;
function slv_to_uint1629_t(x : std_logic_vector) return uint1629_t;
subtype int1629_t is signed(1628 downto 0);
constant int1629_t_SLV_LEN : integer := 1629;
function int1629_t_to_slv(x : int1629_t) return std_logic_vector;
function slv_to_int1629_t(x : std_logic_vector) return int1629_t;
subtype uint1630_t is unsigned(1629 downto 0);
constant uint1630_t_SLV_LEN : integer := 1630;
function uint1630_t_to_slv(x : uint1630_t) return std_logic_vector;
function slv_to_uint1630_t(x : std_logic_vector) return uint1630_t;
subtype int1630_t is signed(1629 downto 0);
constant int1630_t_SLV_LEN : integer := 1630;
function int1630_t_to_slv(x : int1630_t) return std_logic_vector;
function slv_to_int1630_t(x : std_logic_vector) return int1630_t;
subtype uint1631_t is unsigned(1630 downto 0);
constant uint1631_t_SLV_LEN : integer := 1631;
function uint1631_t_to_slv(x : uint1631_t) return std_logic_vector;
function slv_to_uint1631_t(x : std_logic_vector) return uint1631_t;
subtype int1631_t is signed(1630 downto 0);
constant int1631_t_SLV_LEN : integer := 1631;
function int1631_t_to_slv(x : int1631_t) return std_logic_vector;
function slv_to_int1631_t(x : std_logic_vector) return int1631_t;
subtype uint1632_t is unsigned(1631 downto 0);
constant uint1632_t_SLV_LEN : integer := 1632;
function uint1632_t_to_slv(x : uint1632_t) return std_logic_vector;
function slv_to_uint1632_t(x : std_logic_vector) return uint1632_t;
subtype int1632_t is signed(1631 downto 0);
constant int1632_t_SLV_LEN : integer := 1632;
function int1632_t_to_slv(x : int1632_t) return std_logic_vector;
function slv_to_int1632_t(x : std_logic_vector) return int1632_t;
subtype uint1633_t is unsigned(1632 downto 0);
constant uint1633_t_SLV_LEN : integer := 1633;
function uint1633_t_to_slv(x : uint1633_t) return std_logic_vector;
function slv_to_uint1633_t(x : std_logic_vector) return uint1633_t;
subtype int1633_t is signed(1632 downto 0);
constant int1633_t_SLV_LEN : integer := 1633;
function int1633_t_to_slv(x : int1633_t) return std_logic_vector;
function slv_to_int1633_t(x : std_logic_vector) return int1633_t;
subtype uint1634_t is unsigned(1633 downto 0);
constant uint1634_t_SLV_LEN : integer := 1634;
function uint1634_t_to_slv(x : uint1634_t) return std_logic_vector;
function slv_to_uint1634_t(x : std_logic_vector) return uint1634_t;
subtype int1634_t is signed(1633 downto 0);
constant int1634_t_SLV_LEN : integer := 1634;
function int1634_t_to_slv(x : int1634_t) return std_logic_vector;
function slv_to_int1634_t(x : std_logic_vector) return int1634_t;
subtype uint1635_t is unsigned(1634 downto 0);
constant uint1635_t_SLV_LEN : integer := 1635;
function uint1635_t_to_slv(x : uint1635_t) return std_logic_vector;
function slv_to_uint1635_t(x : std_logic_vector) return uint1635_t;
subtype int1635_t is signed(1634 downto 0);
constant int1635_t_SLV_LEN : integer := 1635;
function int1635_t_to_slv(x : int1635_t) return std_logic_vector;
function slv_to_int1635_t(x : std_logic_vector) return int1635_t;
subtype uint1636_t is unsigned(1635 downto 0);
constant uint1636_t_SLV_LEN : integer := 1636;
function uint1636_t_to_slv(x : uint1636_t) return std_logic_vector;
function slv_to_uint1636_t(x : std_logic_vector) return uint1636_t;
subtype int1636_t is signed(1635 downto 0);
constant int1636_t_SLV_LEN : integer := 1636;
function int1636_t_to_slv(x : int1636_t) return std_logic_vector;
function slv_to_int1636_t(x : std_logic_vector) return int1636_t;
subtype uint1637_t is unsigned(1636 downto 0);
constant uint1637_t_SLV_LEN : integer := 1637;
function uint1637_t_to_slv(x : uint1637_t) return std_logic_vector;
function slv_to_uint1637_t(x : std_logic_vector) return uint1637_t;
subtype int1637_t is signed(1636 downto 0);
constant int1637_t_SLV_LEN : integer := 1637;
function int1637_t_to_slv(x : int1637_t) return std_logic_vector;
function slv_to_int1637_t(x : std_logic_vector) return int1637_t;
subtype uint1638_t is unsigned(1637 downto 0);
constant uint1638_t_SLV_LEN : integer := 1638;
function uint1638_t_to_slv(x : uint1638_t) return std_logic_vector;
function slv_to_uint1638_t(x : std_logic_vector) return uint1638_t;
subtype int1638_t is signed(1637 downto 0);
constant int1638_t_SLV_LEN : integer := 1638;
function int1638_t_to_slv(x : int1638_t) return std_logic_vector;
function slv_to_int1638_t(x : std_logic_vector) return int1638_t;
subtype uint1639_t is unsigned(1638 downto 0);
constant uint1639_t_SLV_LEN : integer := 1639;
function uint1639_t_to_slv(x : uint1639_t) return std_logic_vector;
function slv_to_uint1639_t(x : std_logic_vector) return uint1639_t;
subtype int1639_t is signed(1638 downto 0);
constant int1639_t_SLV_LEN : integer := 1639;
function int1639_t_to_slv(x : int1639_t) return std_logic_vector;
function slv_to_int1639_t(x : std_logic_vector) return int1639_t;
subtype uint1640_t is unsigned(1639 downto 0);
constant uint1640_t_SLV_LEN : integer := 1640;
function uint1640_t_to_slv(x : uint1640_t) return std_logic_vector;
function slv_to_uint1640_t(x : std_logic_vector) return uint1640_t;
subtype int1640_t is signed(1639 downto 0);
constant int1640_t_SLV_LEN : integer := 1640;
function int1640_t_to_slv(x : int1640_t) return std_logic_vector;
function slv_to_int1640_t(x : std_logic_vector) return int1640_t;
subtype uint1641_t is unsigned(1640 downto 0);
constant uint1641_t_SLV_LEN : integer := 1641;
function uint1641_t_to_slv(x : uint1641_t) return std_logic_vector;
function slv_to_uint1641_t(x : std_logic_vector) return uint1641_t;
subtype int1641_t is signed(1640 downto 0);
constant int1641_t_SLV_LEN : integer := 1641;
function int1641_t_to_slv(x : int1641_t) return std_logic_vector;
function slv_to_int1641_t(x : std_logic_vector) return int1641_t;
subtype uint1642_t is unsigned(1641 downto 0);
constant uint1642_t_SLV_LEN : integer := 1642;
function uint1642_t_to_slv(x : uint1642_t) return std_logic_vector;
function slv_to_uint1642_t(x : std_logic_vector) return uint1642_t;
subtype int1642_t is signed(1641 downto 0);
constant int1642_t_SLV_LEN : integer := 1642;
function int1642_t_to_slv(x : int1642_t) return std_logic_vector;
function slv_to_int1642_t(x : std_logic_vector) return int1642_t;
subtype uint1643_t is unsigned(1642 downto 0);
constant uint1643_t_SLV_LEN : integer := 1643;
function uint1643_t_to_slv(x : uint1643_t) return std_logic_vector;
function slv_to_uint1643_t(x : std_logic_vector) return uint1643_t;
subtype int1643_t is signed(1642 downto 0);
constant int1643_t_SLV_LEN : integer := 1643;
function int1643_t_to_slv(x : int1643_t) return std_logic_vector;
function slv_to_int1643_t(x : std_logic_vector) return int1643_t;
subtype uint1644_t is unsigned(1643 downto 0);
constant uint1644_t_SLV_LEN : integer := 1644;
function uint1644_t_to_slv(x : uint1644_t) return std_logic_vector;
function slv_to_uint1644_t(x : std_logic_vector) return uint1644_t;
subtype int1644_t is signed(1643 downto 0);
constant int1644_t_SLV_LEN : integer := 1644;
function int1644_t_to_slv(x : int1644_t) return std_logic_vector;
function slv_to_int1644_t(x : std_logic_vector) return int1644_t;
subtype uint1645_t is unsigned(1644 downto 0);
constant uint1645_t_SLV_LEN : integer := 1645;
function uint1645_t_to_slv(x : uint1645_t) return std_logic_vector;
function slv_to_uint1645_t(x : std_logic_vector) return uint1645_t;
subtype int1645_t is signed(1644 downto 0);
constant int1645_t_SLV_LEN : integer := 1645;
function int1645_t_to_slv(x : int1645_t) return std_logic_vector;
function slv_to_int1645_t(x : std_logic_vector) return int1645_t;
subtype uint1646_t is unsigned(1645 downto 0);
constant uint1646_t_SLV_LEN : integer := 1646;
function uint1646_t_to_slv(x : uint1646_t) return std_logic_vector;
function slv_to_uint1646_t(x : std_logic_vector) return uint1646_t;
subtype int1646_t is signed(1645 downto 0);
constant int1646_t_SLV_LEN : integer := 1646;
function int1646_t_to_slv(x : int1646_t) return std_logic_vector;
function slv_to_int1646_t(x : std_logic_vector) return int1646_t;
subtype uint1647_t is unsigned(1646 downto 0);
constant uint1647_t_SLV_LEN : integer := 1647;
function uint1647_t_to_slv(x : uint1647_t) return std_logic_vector;
function slv_to_uint1647_t(x : std_logic_vector) return uint1647_t;
subtype int1647_t is signed(1646 downto 0);
constant int1647_t_SLV_LEN : integer := 1647;
function int1647_t_to_slv(x : int1647_t) return std_logic_vector;
function slv_to_int1647_t(x : std_logic_vector) return int1647_t;
subtype uint1648_t is unsigned(1647 downto 0);
constant uint1648_t_SLV_LEN : integer := 1648;
function uint1648_t_to_slv(x : uint1648_t) return std_logic_vector;
function slv_to_uint1648_t(x : std_logic_vector) return uint1648_t;
subtype int1648_t is signed(1647 downto 0);
constant int1648_t_SLV_LEN : integer := 1648;
function int1648_t_to_slv(x : int1648_t) return std_logic_vector;
function slv_to_int1648_t(x : std_logic_vector) return int1648_t;
subtype uint1649_t is unsigned(1648 downto 0);
constant uint1649_t_SLV_LEN : integer := 1649;
function uint1649_t_to_slv(x : uint1649_t) return std_logic_vector;
function slv_to_uint1649_t(x : std_logic_vector) return uint1649_t;
subtype int1649_t is signed(1648 downto 0);
constant int1649_t_SLV_LEN : integer := 1649;
function int1649_t_to_slv(x : int1649_t) return std_logic_vector;
function slv_to_int1649_t(x : std_logic_vector) return int1649_t;
subtype uint1650_t is unsigned(1649 downto 0);
constant uint1650_t_SLV_LEN : integer := 1650;
function uint1650_t_to_slv(x : uint1650_t) return std_logic_vector;
function slv_to_uint1650_t(x : std_logic_vector) return uint1650_t;
subtype int1650_t is signed(1649 downto 0);
constant int1650_t_SLV_LEN : integer := 1650;
function int1650_t_to_slv(x : int1650_t) return std_logic_vector;
function slv_to_int1650_t(x : std_logic_vector) return int1650_t;
subtype uint1651_t is unsigned(1650 downto 0);
constant uint1651_t_SLV_LEN : integer := 1651;
function uint1651_t_to_slv(x : uint1651_t) return std_logic_vector;
function slv_to_uint1651_t(x : std_logic_vector) return uint1651_t;
subtype int1651_t is signed(1650 downto 0);
constant int1651_t_SLV_LEN : integer := 1651;
function int1651_t_to_slv(x : int1651_t) return std_logic_vector;
function slv_to_int1651_t(x : std_logic_vector) return int1651_t;
subtype uint1652_t is unsigned(1651 downto 0);
constant uint1652_t_SLV_LEN : integer := 1652;
function uint1652_t_to_slv(x : uint1652_t) return std_logic_vector;
function slv_to_uint1652_t(x : std_logic_vector) return uint1652_t;
subtype int1652_t is signed(1651 downto 0);
constant int1652_t_SLV_LEN : integer := 1652;
function int1652_t_to_slv(x : int1652_t) return std_logic_vector;
function slv_to_int1652_t(x : std_logic_vector) return int1652_t;
subtype uint1653_t is unsigned(1652 downto 0);
constant uint1653_t_SLV_LEN : integer := 1653;
function uint1653_t_to_slv(x : uint1653_t) return std_logic_vector;
function slv_to_uint1653_t(x : std_logic_vector) return uint1653_t;
subtype int1653_t is signed(1652 downto 0);
constant int1653_t_SLV_LEN : integer := 1653;
function int1653_t_to_slv(x : int1653_t) return std_logic_vector;
function slv_to_int1653_t(x : std_logic_vector) return int1653_t;
subtype uint1654_t is unsigned(1653 downto 0);
constant uint1654_t_SLV_LEN : integer := 1654;
function uint1654_t_to_slv(x : uint1654_t) return std_logic_vector;
function slv_to_uint1654_t(x : std_logic_vector) return uint1654_t;
subtype int1654_t is signed(1653 downto 0);
constant int1654_t_SLV_LEN : integer := 1654;
function int1654_t_to_slv(x : int1654_t) return std_logic_vector;
function slv_to_int1654_t(x : std_logic_vector) return int1654_t;
subtype uint1655_t is unsigned(1654 downto 0);
constant uint1655_t_SLV_LEN : integer := 1655;
function uint1655_t_to_slv(x : uint1655_t) return std_logic_vector;
function slv_to_uint1655_t(x : std_logic_vector) return uint1655_t;
subtype int1655_t is signed(1654 downto 0);
constant int1655_t_SLV_LEN : integer := 1655;
function int1655_t_to_slv(x : int1655_t) return std_logic_vector;
function slv_to_int1655_t(x : std_logic_vector) return int1655_t;
subtype uint1656_t is unsigned(1655 downto 0);
constant uint1656_t_SLV_LEN : integer := 1656;
function uint1656_t_to_slv(x : uint1656_t) return std_logic_vector;
function slv_to_uint1656_t(x : std_logic_vector) return uint1656_t;
subtype int1656_t is signed(1655 downto 0);
constant int1656_t_SLV_LEN : integer := 1656;
function int1656_t_to_slv(x : int1656_t) return std_logic_vector;
function slv_to_int1656_t(x : std_logic_vector) return int1656_t;
subtype uint1657_t is unsigned(1656 downto 0);
constant uint1657_t_SLV_LEN : integer := 1657;
function uint1657_t_to_slv(x : uint1657_t) return std_logic_vector;
function slv_to_uint1657_t(x : std_logic_vector) return uint1657_t;
subtype int1657_t is signed(1656 downto 0);
constant int1657_t_SLV_LEN : integer := 1657;
function int1657_t_to_slv(x : int1657_t) return std_logic_vector;
function slv_to_int1657_t(x : std_logic_vector) return int1657_t;
subtype uint1658_t is unsigned(1657 downto 0);
constant uint1658_t_SLV_LEN : integer := 1658;
function uint1658_t_to_slv(x : uint1658_t) return std_logic_vector;
function slv_to_uint1658_t(x : std_logic_vector) return uint1658_t;
subtype int1658_t is signed(1657 downto 0);
constant int1658_t_SLV_LEN : integer := 1658;
function int1658_t_to_slv(x : int1658_t) return std_logic_vector;
function slv_to_int1658_t(x : std_logic_vector) return int1658_t;
subtype uint1659_t is unsigned(1658 downto 0);
constant uint1659_t_SLV_LEN : integer := 1659;
function uint1659_t_to_slv(x : uint1659_t) return std_logic_vector;
function slv_to_uint1659_t(x : std_logic_vector) return uint1659_t;
subtype int1659_t is signed(1658 downto 0);
constant int1659_t_SLV_LEN : integer := 1659;
function int1659_t_to_slv(x : int1659_t) return std_logic_vector;
function slv_to_int1659_t(x : std_logic_vector) return int1659_t;
subtype uint1660_t is unsigned(1659 downto 0);
constant uint1660_t_SLV_LEN : integer := 1660;
function uint1660_t_to_slv(x : uint1660_t) return std_logic_vector;
function slv_to_uint1660_t(x : std_logic_vector) return uint1660_t;
subtype int1660_t is signed(1659 downto 0);
constant int1660_t_SLV_LEN : integer := 1660;
function int1660_t_to_slv(x : int1660_t) return std_logic_vector;
function slv_to_int1660_t(x : std_logic_vector) return int1660_t;
subtype uint1661_t is unsigned(1660 downto 0);
constant uint1661_t_SLV_LEN : integer := 1661;
function uint1661_t_to_slv(x : uint1661_t) return std_logic_vector;
function slv_to_uint1661_t(x : std_logic_vector) return uint1661_t;
subtype int1661_t is signed(1660 downto 0);
constant int1661_t_SLV_LEN : integer := 1661;
function int1661_t_to_slv(x : int1661_t) return std_logic_vector;
function slv_to_int1661_t(x : std_logic_vector) return int1661_t;
subtype uint1662_t is unsigned(1661 downto 0);
constant uint1662_t_SLV_LEN : integer := 1662;
function uint1662_t_to_slv(x : uint1662_t) return std_logic_vector;
function slv_to_uint1662_t(x : std_logic_vector) return uint1662_t;
subtype int1662_t is signed(1661 downto 0);
constant int1662_t_SLV_LEN : integer := 1662;
function int1662_t_to_slv(x : int1662_t) return std_logic_vector;
function slv_to_int1662_t(x : std_logic_vector) return int1662_t;
subtype uint1663_t is unsigned(1662 downto 0);
constant uint1663_t_SLV_LEN : integer := 1663;
function uint1663_t_to_slv(x : uint1663_t) return std_logic_vector;
function slv_to_uint1663_t(x : std_logic_vector) return uint1663_t;
subtype int1663_t is signed(1662 downto 0);
constant int1663_t_SLV_LEN : integer := 1663;
function int1663_t_to_slv(x : int1663_t) return std_logic_vector;
function slv_to_int1663_t(x : std_logic_vector) return int1663_t;
subtype uint1664_t is unsigned(1663 downto 0);
constant uint1664_t_SLV_LEN : integer := 1664;
function uint1664_t_to_slv(x : uint1664_t) return std_logic_vector;
function slv_to_uint1664_t(x : std_logic_vector) return uint1664_t;
subtype int1664_t is signed(1663 downto 0);
constant int1664_t_SLV_LEN : integer := 1664;
function int1664_t_to_slv(x : int1664_t) return std_logic_vector;
function slv_to_int1664_t(x : std_logic_vector) return int1664_t;
subtype uint1665_t is unsigned(1664 downto 0);
constant uint1665_t_SLV_LEN : integer := 1665;
function uint1665_t_to_slv(x : uint1665_t) return std_logic_vector;
function slv_to_uint1665_t(x : std_logic_vector) return uint1665_t;
subtype int1665_t is signed(1664 downto 0);
constant int1665_t_SLV_LEN : integer := 1665;
function int1665_t_to_slv(x : int1665_t) return std_logic_vector;
function slv_to_int1665_t(x : std_logic_vector) return int1665_t;
subtype uint1666_t is unsigned(1665 downto 0);
constant uint1666_t_SLV_LEN : integer := 1666;
function uint1666_t_to_slv(x : uint1666_t) return std_logic_vector;
function slv_to_uint1666_t(x : std_logic_vector) return uint1666_t;
subtype int1666_t is signed(1665 downto 0);
constant int1666_t_SLV_LEN : integer := 1666;
function int1666_t_to_slv(x : int1666_t) return std_logic_vector;
function slv_to_int1666_t(x : std_logic_vector) return int1666_t;
subtype uint1667_t is unsigned(1666 downto 0);
constant uint1667_t_SLV_LEN : integer := 1667;
function uint1667_t_to_slv(x : uint1667_t) return std_logic_vector;
function slv_to_uint1667_t(x : std_logic_vector) return uint1667_t;
subtype int1667_t is signed(1666 downto 0);
constant int1667_t_SLV_LEN : integer := 1667;
function int1667_t_to_slv(x : int1667_t) return std_logic_vector;
function slv_to_int1667_t(x : std_logic_vector) return int1667_t;
subtype uint1668_t is unsigned(1667 downto 0);
constant uint1668_t_SLV_LEN : integer := 1668;
function uint1668_t_to_slv(x : uint1668_t) return std_logic_vector;
function slv_to_uint1668_t(x : std_logic_vector) return uint1668_t;
subtype int1668_t is signed(1667 downto 0);
constant int1668_t_SLV_LEN : integer := 1668;
function int1668_t_to_slv(x : int1668_t) return std_logic_vector;
function slv_to_int1668_t(x : std_logic_vector) return int1668_t;
subtype uint1669_t is unsigned(1668 downto 0);
constant uint1669_t_SLV_LEN : integer := 1669;
function uint1669_t_to_slv(x : uint1669_t) return std_logic_vector;
function slv_to_uint1669_t(x : std_logic_vector) return uint1669_t;
subtype int1669_t is signed(1668 downto 0);
constant int1669_t_SLV_LEN : integer := 1669;
function int1669_t_to_slv(x : int1669_t) return std_logic_vector;
function slv_to_int1669_t(x : std_logic_vector) return int1669_t;
subtype uint1670_t is unsigned(1669 downto 0);
constant uint1670_t_SLV_LEN : integer := 1670;
function uint1670_t_to_slv(x : uint1670_t) return std_logic_vector;
function slv_to_uint1670_t(x : std_logic_vector) return uint1670_t;
subtype int1670_t is signed(1669 downto 0);
constant int1670_t_SLV_LEN : integer := 1670;
function int1670_t_to_slv(x : int1670_t) return std_logic_vector;
function slv_to_int1670_t(x : std_logic_vector) return int1670_t;
subtype uint1671_t is unsigned(1670 downto 0);
constant uint1671_t_SLV_LEN : integer := 1671;
function uint1671_t_to_slv(x : uint1671_t) return std_logic_vector;
function slv_to_uint1671_t(x : std_logic_vector) return uint1671_t;
subtype int1671_t is signed(1670 downto 0);
constant int1671_t_SLV_LEN : integer := 1671;
function int1671_t_to_slv(x : int1671_t) return std_logic_vector;
function slv_to_int1671_t(x : std_logic_vector) return int1671_t;
subtype uint1672_t is unsigned(1671 downto 0);
constant uint1672_t_SLV_LEN : integer := 1672;
function uint1672_t_to_slv(x : uint1672_t) return std_logic_vector;
function slv_to_uint1672_t(x : std_logic_vector) return uint1672_t;
subtype int1672_t is signed(1671 downto 0);
constant int1672_t_SLV_LEN : integer := 1672;
function int1672_t_to_slv(x : int1672_t) return std_logic_vector;
function slv_to_int1672_t(x : std_logic_vector) return int1672_t;
subtype uint1673_t is unsigned(1672 downto 0);
constant uint1673_t_SLV_LEN : integer := 1673;
function uint1673_t_to_slv(x : uint1673_t) return std_logic_vector;
function slv_to_uint1673_t(x : std_logic_vector) return uint1673_t;
subtype int1673_t is signed(1672 downto 0);
constant int1673_t_SLV_LEN : integer := 1673;
function int1673_t_to_slv(x : int1673_t) return std_logic_vector;
function slv_to_int1673_t(x : std_logic_vector) return int1673_t;
subtype uint1674_t is unsigned(1673 downto 0);
constant uint1674_t_SLV_LEN : integer := 1674;
function uint1674_t_to_slv(x : uint1674_t) return std_logic_vector;
function slv_to_uint1674_t(x : std_logic_vector) return uint1674_t;
subtype int1674_t is signed(1673 downto 0);
constant int1674_t_SLV_LEN : integer := 1674;
function int1674_t_to_slv(x : int1674_t) return std_logic_vector;
function slv_to_int1674_t(x : std_logic_vector) return int1674_t;
subtype uint1675_t is unsigned(1674 downto 0);
constant uint1675_t_SLV_LEN : integer := 1675;
function uint1675_t_to_slv(x : uint1675_t) return std_logic_vector;
function slv_to_uint1675_t(x : std_logic_vector) return uint1675_t;
subtype int1675_t is signed(1674 downto 0);
constant int1675_t_SLV_LEN : integer := 1675;
function int1675_t_to_slv(x : int1675_t) return std_logic_vector;
function slv_to_int1675_t(x : std_logic_vector) return int1675_t;
subtype uint1676_t is unsigned(1675 downto 0);
constant uint1676_t_SLV_LEN : integer := 1676;
function uint1676_t_to_slv(x : uint1676_t) return std_logic_vector;
function slv_to_uint1676_t(x : std_logic_vector) return uint1676_t;
subtype int1676_t is signed(1675 downto 0);
constant int1676_t_SLV_LEN : integer := 1676;
function int1676_t_to_slv(x : int1676_t) return std_logic_vector;
function slv_to_int1676_t(x : std_logic_vector) return int1676_t;
subtype uint1677_t is unsigned(1676 downto 0);
constant uint1677_t_SLV_LEN : integer := 1677;
function uint1677_t_to_slv(x : uint1677_t) return std_logic_vector;
function slv_to_uint1677_t(x : std_logic_vector) return uint1677_t;
subtype int1677_t is signed(1676 downto 0);
constant int1677_t_SLV_LEN : integer := 1677;
function int1677_t_to_slv(x : int1677_t) return std_logic_vector;
function slv_to_int1677_t(x : std_logic_vector) return int1677_t;
subtype uint1678_t is unsigned(1677 downto 0);
constant uint1678_t_SLV_LEN : integer := 1678;
function uint1678_t_to_slv(x : uint1678_t) return std_logic_vector;
function slv_to_uint1678_t(x : std_logic_vector) return uint1678_t;
subtype int1678_t is signed(1677 downto 0);
constant int1678_t_SLV_LEN : integer := 1678;
function int1678_t_to_slv(x : int1678_t) return std_logic_vector;
function slv_to_int1678_t(x : std_logic_vector) return int1678_t;
subtype uint1679_t is unsigned(1678 downto 0);
constant uint1679_t_SLV_LEN : integer := 1679;
function uint1679_t_to_slv(x : uint1679_t) return std_logic_vector;
function slv_to_uint1679_t(x : std_logic_vector) return uint1679_t;
subtype int1679_t is signed(1678 downto 0);
constant int1679_t_SLV_LEN : integer := 1679;
function int1679_t_to_slv(x : int1679_t) return std_logic_vector;
function slv_to_int1679_t(x : std_logic_vector) return int1679_t;
subtype uint1680_t is unsigned(1679 downto 0);
constant uint1680_t_SLV_LEN : integer := 1680;
function uint1680_t_to_slv(x : uint1680_t) return std_logic_vector;
function slv_to_uint1680_t(x : std_logic_vector) return uint1680_t;
subtype int1680_t is signed(1679 downto 0);
constant int1680_t_SLV_LEN : integer := 1680;
function int1680_t_to_slv(x : int1680_t) return std_logic_vector;
function slv_to_int1680_t(x : std_logic_vector) return int1680_t;
subtype uint1681_t is unsigned(1680 downto 0);
constant uint1681_t_SLV_LEN : integer := 1681;
function uint1681_t_to_slv(x : uint1681_t) return std_logic_vector;
function slv_to_uint1681_t(x : std_logic_vector) return uint1681_t;
subtype int1681_t is signed(1680 downto 0);
constant int1681_t_SLV_LEN : integer := 1681;
function int1681_t_to_slv(x : int1681_t) return std_logic_vector;
function slv_to_int1681_t(x : std_logic_vector) return int1681_t;
subtype uint1682_t is unsigned(1681 downto 0);
constant uint1682_t_SLV_LEN : integer := 1682;
function uint1682_t_to_slv(x : uint1682_t) return std_logic_vector;
function slv_to_uint1682_t(x : std_logic_vector) return uint1682_t;
subtype int1682_t is signed(1681 downto 0);
constant int1682_t_SLV_LEN : integer := 1682;
function int1682_t_to_slv(x : int1682_t) return std_logic_vector;
function slv_to_int1682_t(x : std_logic_vector) return int1682_t;
subtype uint1683_t is unsigned(1682 downto 0);
constant uint1683_t_SLV_LEN : integer := 1683;
function uint1683_t_to_slv(x : uint1683_t) return std_logic_vector;
function slv_to_uint1683_t(x : std_logic_vector) return uint1683_t;
subtype int1683_t is signed(1682 downto 0);
constant int1683_t_SLV_LEN : integer := 1683;
function int1683_t_to_slv(x : int1683_t) return std_logic_vector;
function slv_to_int1683_t(x : std_logic_vector) return int1683_t;
subtype uint1684_t is unsigned(1683 downto 0);
constant uint1684_t_SLV_LEN : integer := 1684;
function uint1684_t_to_slv(x : uint1684_t) return std_logic_vector;
function slv_to_uint1684_t(x : std_logic_vector) return uint1684_t;
subtype int1684_t is signed(1683 downto 0);
constant int1684_t_SLV_LEN : integer := 1684;
function int1684_t_to_slv(x : int1684_t) return std_logic_vector;
function slv_to_int1684_t(x : std_logic_vector) return int1684_t;
subtype uint1685_t is unsigned(1684 downto 0);
constant uint1685_t_SLV_LEN : integer := 1685;
function uint1685_t_to_slv(x : uint1685_t) return std_logic_vector;
function slv_to_uint1685_t(x : std_logic_vector) return uint1685_t;
subtype int1685_t is signed(1684 downto 0);
constant int1685_t_SLV_LEN : integer := 1685;
function int1685_t_to_slv(x : int1685_t) return std_logic_vector;
function slv_to_int1685_t(x : std_logic_vector) return int1685_t;
subtype uint1686_t is unsigned(1685 downto 0);
constant uint1686_t_SLV_LEN : integer := 1686;
function uint1686_t_to_slv(x : uint1686_t) return std_logic_vector;
function slv_to_uint1686_t(x : std_logic_vector) return uint1686_t;
subtype int1686_t is signed(1685 downto 0);
constant int1686_t_SLV_LEN : integer := 1686;
function int1686_t_to_slv(x : int1686_t) return std_logic_vector;
function slv_to_int1686_t(x : std_logic_vector) return int1686_t;
subtype uint1687_t is unsigned(1686 downto 0);
constant uint1687_t_SLV_LEN : integer := 1687;
function uint1687_t_to_slv(x : uint1687_t) return std_logic_vector;
function slv_to_uint1687_t(x : std_logic_vector) return uint1687_t;
subtype int1687_t is signed(1686 downto 0);
constant int1687_t_SLV_LEN : integer := 1687;
function int1687_t_to_slv(x : int1687_t) return std_logic_vector;
function slv_to_int1687_t(x : std_logic_vector) return int1687_t;
subtype uint1688_t is unsigned(1687 downto 0);
constant uint1688_t_SLV_LEN : integer := 1688;
function uint1688_t_to_slv(x : uint1688_t) return std_logic_vector;
function slv_to_uint1688_t(x : std_logic_vector) return uint1688_t;
subtype int1688_t is signed(1687 downto 0);
constant int1688_t_SLV_LEN : integer := 1688;
function int1688_t_to_slv(x : int1688_t) return std_logic_vector;
function slv_to_int1688_t(x : std_logic_vector) return int1688_t;
subtype uint1689_t is unsigned(1688 downto 0);
constant uint1689_t_SLV_LEN : integer := 1689;
function uint1689_t_to_slv(x : uint1689_t) return std_logic_vector;
function slv_to_uint1689_t(x : std_logic_vector) return uint1689_t;
subtype int1689_t is signed(1688 downto 0);
constant int1689_t_SLV_LEN : integer := 1689;
function int1689_t_to_slv(x : int1689_t) return std_logic_vector;
function slv_to_int1689_t(x : std_logic_vector) return int1689_t;
subtype uint1690_t is unsigned(1689 downto 0);
constant uint1690_t_SLV_LEN : integer := 1690;
function uint1690_t_to_slv(x : uint1690_t) return std_logic_vector;
function slv_to_uint1690_t(x : std_logic_vector) return uint1690_t;
subtype int1690_t is signed(1689 downto 0);
constant int1690_t_SLV_LEN : integer := 1690;
function int1690_t_to_slv(x : int1690_t) return std_logic_vector;
function slv_to_int1690_t(x : std_logic_vector) return int1690_t;
subtype uint1691_t is unsigned(1690 downto 0);
constant uint1691_t_SLV_LEN : integer := 1691;
function uint1691_t_to_slv(x : uint1691_t) return std_logic_vector;
function slv_to_uint1691_t(x : std_logic_vector) return uint1691_t;
subtype int1691_t is signed(1690 downto 0);
constant int1691_t_SLV_LEN : integer := 1691;
function int1691_t_to_slv(x : int1691_t) return std_logic_vector;
function slv_to_int1691_t(x : std_logic_vector) return int1691_t;
subtype uint1692_t is unsigned(1691 downto 0);
constant uint1692_t_SLV_LEN : integer := 1692;
function uint1692_t_to_slv(x : uint1692_t) return std_logic_vector;
function slv_to_uint1692_t(x : std_logic_vector) return uint1692_t;
subtype int1692_t is signed(1691 downto 0);
constant int1692_t_SLV_LEN : integer := 1692;
function int1692_t_to_slv(x : int1692_t) return std_logic_vector;
function slv_to_int1692_t(x : std_logic_vector) return int1692_t;
subtype uint1693_t is unsigned(1692 downto 0);
constant uint1693_t_SLV_LEN : integer := 1693;
function uint1693_t_to_slv(x : uint1693_t) return std_logic_vector;
function slv_to_uint1693_t(x : std_logic_vector) return uint1693_t;
subtype int1693_t is signed(1692 downto 0);
constant int1693_t_SLV_LEN : integer := 1693;
function int1693_t_to_slv(x : int1693_t) return std_logic_vector;
function slv_to_int1693_t(x : std_logic_vector) return int1693_t;
subtype uint1694_t is unsigned(1693 downto 0);
constant uint1694_t_SLV_LEN : integer := 1694;
function uint1694_t_to_slv(x : uint1694_t) return std_logic_vector;
function slv_to_uint1694_t(x : std_logic_vector) return uint1694_t;
subtype int1694_t is signed(1693 downto 0);
constant int1694_t_SLV_LEN : integer := 1694;
function int1694_t_to_slv(x : int1694_t) return std_logic_vector;
function slv_to_int1694_t(x : std_logic_vector) return int1694_t;
subtype uint1695_t is unsigned(1694 downto 0);
constant uint1695_t_SLV_LEN : integer := 1695;
function uint1695_t_to_slv(x : uint1695_t) return std_logic_vector;
function slv_to_uint1695_t(x : std_logic_vector) return uint1695_t;
subtype int1695_t is signed(1694 downto 0);
constant int1695_t_SLV_LEN : integer := 1695;
function int1695_t_to_slv(x : int1695_t) return std_logic_vector;
function slv_to_int1695_t(x : std_logic_vector) return int1695_t;
subtype uint1696_t is unsigned(1695 downto 0);
constant uint1696_t_SLV_LEN : integer := 1696;
function uint1696_t_to_slv(x : uint1696_t) return std_logic_vector;
function slv_to_uint1696_t(x : std_logic_vector) return uint1696_t;
subtype int1696_t is signed(1695 downto 0);
constant int1696_t_SLV_LEN : integer := 1696;
function int1696_t_to_slv(x : int1696_t) return std_logic_vector;
function slv_to_int1696_t(x : std_logic_vector) return int1696_t;
subtype uint1697_t is unsigned(1696 downto 0);
constant uint1697_t_SLV_LEN : integer := 1697;
function uint1697_t_to_slv(x : uint1697_t) return std_logic_vector;
function slv_to_uint1697_t(x : std_logic_vector) return uint1697_t;
subtype int1697_t is signed(1696 downto 0);
constant int1697_t_SLV_LEN : integer := 1697;
function int1697_t_to_slv(x : int1697_t) return std_logic_vector;
function slv_to_int1697_t(x : std_logic_vector) return int1697_t;
subtype uint1698_t is unsigned(1697 downto 0);
constant uint1698_t_SLV_LEN : integer := 1698;
function uint1698_t_to_slv(x : uint1698_t) return std_logic_vector;
function slv_to_uint1698_t(x : std_logic_vector) return uint1698_t;
subtype int1698_t is signed(1697 downto 0);
constant int1698_t_SLV_LEN : integer := 1698;
function int1698_t_to_slv(x : int1698_t) return std_logic_vector;
function slv_to_int1698_t(x : std_logic_vector) return int1698_t;
subtype uint1699_t is unsigned(1698 downto 0);
constant uint1699_t_SLV_LEN : integer := 1699;
function uint1699_t_to_slv(x : uint1699_t) return std_logic_vector;
function slv_to_uint1699_t(x : std_logic_vector) return uint1699_t;
subtype int1699_t is signed(1698 downto 0);
constant int1699_t_SLV_LEN : integer := 1699;
function int1699_t_to_slv(x : int1699_t) return std_logic_vector;
function slv_to_int1699_t(x : std_logic_vector) return int1699_t;
subtype uint1700_t is unsigned(1699 downto 0);
constant uint1700_t_SLV_LEN : integer := 1700;
function uint1700_t_to_slv(x : uint1700_t) return std_logic_vector;
function slv_to_uint1700_t(x : std_logic_vector) return uint1700_t;
subtype int1700_t is signed(1699 downto 0);
constant int1700_t_SLV_LEN : integer := 1700;
function int1700_t_to_slv(x : int1700_t) return std_logic_vector;
function slv_to_int1700_t(x : std_logic_vector) return int1700_t;
subtype uint1701_t is unsigned(1700 downto 0);
constant uint1701_t_SLV_LEN : integer := 1701;
function uint1701_t_to_slv(x : uint1701_t) return std_logic_vector;
function slv_to_uint1701_t(x : std_logic_vector) return uint1701_t;
subtype int1701_t is signed(1700 downto 0);
constant int1701_t_SLV_LEN : integer := 1701;
function int1701_t_to_slv(x : int1701_t) return std_logic_vector;
function slv_to_int1701_t(x : std_logic_vector) return int1701_t;
subtype uint1702_t is unsigned(1701 downto 0);
constant uint1702_t_SLV_LEN : integer := 1702;
function uint1702_t_to_slv(x : uint1702_t) return std_logic_vector;
function slv_to_uint1702_t(x : std_logic_vector) return uint1702_t;
subtype int1702_t is signed(1701 downto 0);
constant int1702_t_SLV_LEN : integer := 1702;
function int1702_t_to_slv(x : int1702_t) return std_logic_vector;
function slv_to_int1702_t(x : std_logic_vector) return int1702_t;
subtype uint1703_t is unsigned(1702 downto 0);
constant uint1703_t_SLV_LEN : integer := 1703;
function uint1703_t_to_slv(x : uint1703_t) return std_logic_vector;
function slv_to_uint1703_t(x : std_logic_vector) return uint1703_t;
subtype int1703_t is signed(1702 downto 0);
constant int1703_t_SLV_LEN : integer := 1703;
function int1703_t_to_slv(x : int1703_t) return std_logic_vector;
function slv_to_int1703_t(x : std_logic_vector) return int1703_t;
subtype uint1704_t is unsigned(1703 downto 0);
constant uint1704_t_SLV_LEN : integer := 1704;
function uint1704_t_to_slv(x : uint1704_t) return std_logic_vector;
function slv_to_uint1704_t(x : std_logic_vector) return uint1704_t;
subtype int1704_t is signed(1703 downto 0);
constant int1704_t_SLV_LEN : integer := 1704;
function int1704_t_to_slv(x : int1704_t) return std_logic_vector;
function slv_to_int1704_t(x : std_logic_vector) return int1704_t;
subtype uint1705_t is unsigned(1704 downto 0);
constant uint1705_t_SLV_LEN : integer := 1705;
function uint1705_t_to_slv(x : uint1705_t) return std_logic_vector;
function slv_to_uint1705_t(x : std_logic_vector) return uint1705_t;
subtype int1705_t is signed(1704 downto 0);
constant int1705_t_SLV_LEN : integer := 1705;
function int1705_t_to_slv(x : int1705_t) return std_logic_vector;
function slv_to_int1705_t(x : std_logic_vector) return int1705_t;
subtype uint1706_t is unsigned(1705 downto 0);
constant uint1706_t_SLV_LEN : integer := 1706;
function uint1706_t_to_slv(x : uint1706_t) return std_logic_vector;
function slv_to_uint1706_t(x : std_logic_vector) return uint1706_t;
subtype int1706_t is signed(1705 downto 0);
constant int1706_t_SLV_LEN : integer := 1706;
function int1706_t_to_slv(x : int1706_t) return std_logic_vector;
function slv_to_int1706_t(x : std_logic_vector) return int1706_t;
subtype uint1707_t is unsigned(1706 downto 0);
constant uint1707_t_SLV_LEN : integer := 1707;
function uint1707_t_to_slv(x : uint1707_t) return std_logic_vector;
function slv_to_uint1707_t(x : std_logic_vector) return uint1707_t;
subtype int1707_t is signed(1706 downto 0);
constant int1707_t_SLV_LEN : integer := 1707;
function int1707_t_to_slv(x : int1707_t) return std_logic_vector;
function slv_to_int1707_t(x : std_logic_vector) return int1707_t;
subtype uint1708_t is unsigned(1707 downto 0);
constant uint1708_t_SLV_LEN : integer := 1708;
function uint1708_t_to_slv(x : uint1708_t) return std_logic_vector;
function slv_to_uint1708_t(x : std_logic_vector) return uint1708_t;
subtype int1708_t is signed(1707 downto 0);
constant int1708_t_SLV_LEN : integer := 1708;
function int1708_t_to_slv(x : int1708_t) return std_logic_vector;
function slv_to_int1708_t(x : std_logic_vector) return int1708_t;
subtype uint1709_t is unsigned(1708 downto 0);
constant uint1709_t_SLV_LEN : integer := 1709;
function uint1709_t_to_slv(x : uint1709_t) return std_logic_vector;
function slv_to_uint1709_t(x : std_logic_vector) return uint1709_t;
subtype int1709_t is signed(1708 downto 0);
constant int1709_t_SLV_LEN : integer := 1709;
function int1709_t_to_slv(x : int1709_t) return std_logic_vector;
function slv_to_int1709_t(x : std_logic_vector) return int1709_t;
subtype uint1710_t is unsigned(1709 downto 0);
constant uint1710_t_SLV_LEN : integer := 1710;
function uint1710_t_to_slv(x : uint1710_t) return std_logic_vector;
function slv_to_uint1710_t(x : std_logic_vector) return uint1710_t;
subtype int1710_t is signed(1709 downto 0);
constant int1710_t_SLV_LEN : integer := 1710;
function int1710_t_to_slv(x : int1710_t) return std_logic_vector;
function slv_to_int1710_t(x : std_logic_vector) return int1710_t;
subtype uint1711_t is unsigned(1710 downto 0);
constant uint1711_t_SLV_LEN : integer := 1711;
function uint1711_t_to_slv(x : uint1711_t) return std_logic_vector;
function slv_to_uint1711_t(x : std_logic_vector) return uint1711_t;
subtype int1711_t is signed(1710 downto 0);
constant int1711_t_SLV_LEN : integer := 1711;
function int1711_t_to_slv(x : int1711_t) return std_logic_vector;
function slv_to_int1711_t(x : std_logic_vector) return int1711_t;
subtype uint1712_t is unsigned(1711 downto 0);
constant uint1712_t_SLV_LEN : integer := 1712;
function uint1712_t_to_slv(x : uint1712_t) return std_logic_vector;
function slv_to_uint1712_t(x : std_logic_vector) return uint1712_t;
subtype int1712_t is signed(1711 downto 0);
constant int1712_t_SLV_LEN : integer := 1712;
function int1712_t_to_slv(x : int1712_t) return std_logic_vector;
function slv_to_int1712_t(x : std_logic_vector) return int1712_t;
subtype uint1713_t is unsigned(1712 downto 0);
constant uint1713_t_SLV_LEN : integer := 1713;
function uint1713_t_to_slv(x : uint1713_t) return std_logic_vector;
function slv_to_uint1713_t(x : std_logic_vector) return uint1713_t;
subtype int1713_t is signed(1712 downto 0);
constant int1713_t_SLV_LEN : integer := 1713;
function int1713_t_to_slv(x : int1713_t) return std_logic_vector;
function slv_to_int1713_t(x : std_logic_vector) return int1713_t;
subtype uint1714_t is unsigned(1713 downto 0);
constant uint1714_t_SLV_LEN : integer := 1714;
function uint1714_t_to_slv(x : uint1714_t) return std_logic_vector;
function slv_to_uint1714_t(x : std_logic_vector) return uint1714_t;
subtype int1714_t is signed(1713 downto 0);
constant int1714_t_SLV_LEN : integer := 1714;
function int1714_t_to_slv(x : int1714_t) return std_logic_vector;
function slv_to_int1714_t(x : std_logic_vector) return int1714_t;
subtype uint1715_t is unsigned(1714 downto 0);
constant uint1715_t_SLV_LEN : integer := 1715;
function uint1715_t_to_slv(x : uint1715_t) return std_logic_vector;
function slv_to_uint1715_t(x : std_logic_vector) return uint1715_t;
subtype int1715_t is signed(1714 downto 0);
constant int1715_t_SLV_LEN : integer := 1715;
function int1715_t_to_slv(x : int1715_t) return std_logic_vector;
function slv_to_int1715_t(x : std_logic_vector) return int1715_t;
subtype uint1716_t is unsigned(1715 downto 0);
constant uint1716_t_SLV_LEN : integer := 1716;
function uint1716_t_to_slv(x : uint1716_t) return std_logic_vector;
function slv_to_uint1716_t(x : std_logic_vector) return uint1716_t;
subtype int1716_t is signed(1715 downto 0);
constant int1716_t_SLV_LEN : integer := 1716;
function int1716_t_to_slv(x : int1716_t) return std_logic_vector;
function slv_to_int1716_t(x : std_logic_vector) return int1716_t;
subtype uint1717_t is unsigned(1716 downto 0);
constant uint1717_t_SLV_LEN : integer := 1717;
function uint1717_t_to_slv(x : uint1717_t) return std_logic_vector;
function slv_to_uint1717_t(x : std_logic_vector) return uint1717_t;
subtype int1717_t is signed(1716 downto 0);
constant int1717_t_SLV_LEN : integer := 1717;
function int1717_t_to_slv(x : int1717_t) return std_logic_vector;
function slv_to_int1717_t(x : std_logic_vector) return int1717_t;
subtype uint1718_t is unsigned(1717 downto 0);
constant uint1718_t_SLV_LEN : integer := 1718;
function uint1718_t_to_slv(x : uint1718_t) return std_logic_vector;
function slv_to_uint1718_t(x : std_logic_vector) return uint1718_t;
subtype int1718_t is signed(1717 downto 0);
constant int1718_t_SLV_LEN : integer := 1718;
function int1718_t_to_slv(x : int1718_t) return std_logic_vector;
function slv_to_int1718_t(x : std_logic_vector) return int1718_t;
subtype uint1719_t is unsigned(1718 downto 0);
constant uint1719_t_SLV_LEN : integer := 1719;
function uint1719_t_to_slv(x : uint1719_t) return std_logic_vector;
function slv_to_uint1719_t(x : std_logic_vector) return uint1719_t;
subtype int1719_t is signed(1718 downto 0);
constant int1719_t_SLV_LEN : integer := 1719;
function int1719_t_to_slv(x : int1719_t) return std_logic_vector;
function slv_to_int1719_t(x : std_logic_vector) return int1719_t;
subtype uint1720_t is unsigned(1719 downto 0);
constant uint1720_t_SLV_LEN : integer := 1720;
function uint1720_t_to_slv(x : uint1720_t) return std_logic_vector;
function slv_to_uint1720_t(x : std_logic_vector) return uint1720_t;
subtype int1720_t is signed(1719 downto 0);
constant int1720_t_SLV_LEN : integer := 1720;
function int1720_t_to_slv(x : int1720_t) return std_logic_vector;
function slv_to_int1720_t(x : std_logic_vector) return int1720_t;
subtype uint1721_t is unsigned(1720 downto 0);
constant uint1721_t_SLV_LEN : integer := 1721;
function uint1721_t_to_slv(x : uint1721_t) return std_logic_vector;
function slv_to_uint1721_t(x : std_logic_vector) return uint1721_t;
subtype int1721_t is signed(1720 downto 0);
constant int1721_t_SLV_LEN : integer := 1721;
function int1721_t_to_slv(x : int1721_t) return std_logic_vector;
function slv_to_int1721_t(x : std_logic_vector) return int1721_t;
subtype uint1722_t is unsigned(1721 downto 0);
constant uint1722_t_SLV_LEN : integer := 1722;
function uint1722_t_to_slv(x : uint1722_t) return std_logic_vector;
function slv_to_uint1722_t(x : std_logic_vector) return uint1722_t;
subtype int1722_t is signed(1721 downto 0);
constant int1722_t_SLV_LEN : integer := 1722;
function int1722_t_to_slv(x : int1722_t) return std_logic_vector;
function slv_to_int1722_t(x : std_logic_vector) return int1722_t;
subtype uint1723_t is unsigned(1722 downto 0);
constant uint1723_t_SLV_LEN : integer := 1723;
function uint1723_t_to_slv(x : uint1723_t) return std_logic_vector;
function slv_to_uint1723_t(x : std_logic_vector) return uint1723_t;
subtype int1723_t is signed(1722 downto 0);
constant int1723_t_SLV_LEN : integer := 1723;
function int1723_t_to_slv(x : int1723_t) return std_logic_vector;
function slv_to_int1723_t(x : std_logic_vector) return int1723_t;
subtype uint1724_t is unsigned(1723 downto 0);
constant uint1724_t_SLV_LEN : integer := 1724;
function uint1724_t_to_slv(x : uint1724_t) return std_logic_vector;
function slv_to_uint1724_t(x : std_logic_vector) return uint1724_t;
subtype int1724_t is signed(1723 downto 0);
constant int1724_t_SLV_LEN : integer := 1724;
function int1724_t_to_slv(x : int1724_t) return std_logic_vector;
function slv_to_int1724_t(x : std_logic_vector) return int1724_t;
subtype uint1725_t is unsigned(1724 downto 0);
constant uint1725_t_SLV_LEN : integer := 1725;
function uint1725_t_to_slv(x : uint1725_t) return std_logic_vector;
function slv_to_uint1725_t(x : std_logic_vector) return uint1725_t;
subtype int1725_t is signed(1724 downto 0);
constant int1725_t_SLV_LEN : integer := 1725;
function int1725_t_to_slv(x : int1725_t) return std_logic_vector;
function slv_to_int1725_t(x : std_logic_vector) return int1725_t;
subtype uint1726_t is unsigned(1725 downto 0);
constant uint1726_t_SLV_LEN : integer := 1726;
function uint1726_t_to_slv(x : uint1726_t) return std_logic_vector;
function slv_to_uint1726_t(x : std_logic_vector) return uint1726_t;
subtype int1726_t is signed(1725 downto 0);
constant int1726_t_SLV_LEN : integer := 1726;
function int1726_t_to_slv(x : int1726_t) return std_logic_vector;
function slv_to_int1726_t(x : std_logic_vector) return int1726_t;
subtype uint1727_t is unsigned(1726 downto 0);
constant uint1727_t_SLV_LEN : integer := 1727;
function uint1727_t_to_slv(x : uint1727_t) return std_logic_vector;
function slv_to_uint1727_t(x : std_logic_vector) return uint1727_t;
subtype int1727_t is signed(1726 downto 0);
constant int1727_t_SLV_LEN : integer := 1727;
function int1727_t_to_slv(x : int1727_t) return std_logic_vector;
function slv_to_int1727_t(x : std_logic_vector) return int1727_t;
subtype uint1728_t is unsigned(1727 downto 0);
constant uint1728_t_SLV_LEN : integer := 1728;
function uint1728_t_to_slv(x : uint1728_t) return std_logic_vector;
function slv_to_uint1728_t(x : std_logic_vector) return uint1728_t;
subtype int1728_t is signed(1727 downto 0);
constant int1728_t_SLV_LEN : integer := 1728;
function int1728_t_to_slv(x : int1728_t) return std_logic_vector;
function slv_to_int1728_t(x : std_logic_vector) return int1728_t;
subtype uint1729_t is unsigned(1728 downto 0);
constant uint1729_t_SLV_LEN : integer := 1729;
function uint1729_t_to_slv(x : uint1729_t) return std_logic_vector;
function slv_to_uint1729_t(x : std_logic_vector) return uint1729_t;
subtype int1729_t is signed(1728 downto 0);
constant int1729_t_SLV_LEN : integer := 1729;
function int1729_t_to_slv(x : int1729_t) return std_logic_vector;
function slv_to_int1729_t(x : std_logic_vector) return int1729_t;
subtype uint1730_t is unsigned(1729 downto 0);
constant uint1730_t_SLV_LEN : integer := 1730;
function uint1730_t_to_slv(x : uint1730_t) return std_logic_vector;
function slv_to_uint1730_t(x : std_logic_vector) return uint1730_t;
subtype int1730_t is signed(1729 downto 0);
constant int1730_t_SLV_LEN : integer := 1730;
function int1730_t_to_slv(x : int1730_t) return std_logic_vector;
function slv_to_int1730_t(x : std_logic_vector) return int1730_t;
subtype uint1731_t is unsigned(1730 downto 0);
constant uint1731_t_SLV_LEN : integer := 1731;
function uint1731_t_to_slv(x : uint1731_t) return std_logic_vector;
function slv_to_uint1731_t(x : std_logic_vector) return uint1731_t;
subtype int1731_t is signed(1730 downto 0);
constant int1731_t_SLV_LEN : integer := 1731;
function int1731_t_to_slv(x : int1731_t) return std_logic_vector;
function slv_to_int1731_t(x : std_logic_vector) return int1731_t;
subtype uint1732_t is unsigned(1731 downto 0);
constant uint1732_t_SLV_LEN : integer := 1732;
function uint1732_t_to_slv(x : uint1732_t) return std_logic_vector;
function slv_to_uint1732_t(x : std_logic_vector) return uint1732_t;
subtype int1732_t is signed(1731 downto 0);
constant int1732_t_SLV_LEN : integer := 1732;
function int1732_t_to_slv(x : int1732_t) return std_logic_vector;
function slv_to_int1732_t(x : std_logic_vector) return int1732_t;
subtype uint1733_t is unsigned(1732 downto 0);
constant uint1733_t_SLV_LEN : integer := 1733;
function uint1733_t_to_slv(x : uint1733_t) return std_logic_vector;
function slv_to_uint1733_t(x : std_logic_vector) return uint1733_t;
subtype int1733_t is signed(1732 downto 0);
constant int1733_t_SLV_LEN : integer := 1733;
function int1733_t_to_slv(x : int1733_t) return std_logic_vector;
function slv_to_int1733_t(x : std_logic_vector) return int1733_t;
subtype uint1734_t is unsigned(1733 downto 0);
constant uint1734_t_SLV_LEN : integer := 1734;
function uint1734_t_to_slv(x : uint1734_t) return std_logic_vector;
function slv_to_uint1734_t(x : std_logic_vector) return uint1734_t;
subtype int1734_t is signed(1733 downto 0);
constant int1734_t_SLV_LEN : integer := 1734;
function int1734_t_to_slv(x : int1734_t) return std_logic_vector;
function slv_to_int1734_t(x : std_logic_vector) return int1734_t;
subtype uint1735_t is unsigned(1734 downto 0);
constant uint1735_t_SLV_LEN : integer := 1735;
function uint1735_t_to_slv(x : uint1735_t) return std_logic_vector;
function slv_to_uint1735_t(x : std_logic_vector) return uint1735_t;
subtype int1735_t is signed(1734 downto 0);
constant int1735_t_SLV_LEN : integer := 1735;
function int1735_t_to_slv(x : int1735_t) return std_logic_vector;
function slv_to_int1735_t(x : std_logic_vector) return int1735_t;
subtype uint1736_t is unsigned(1735 downto 0);
constant uint1736_t_SLV_LEN : integer := 1736;
function uint1736_t_to_slv(x : uint1736_t) return std_logic_vector;
function slv_to_uint1736_t(x : std_logic_vector) return uint1736_t;
subtype int1736_t is signed(1735 downto 0);
constant int1736_t_SLV_LEN : integer := 1736;
function int1736_t_to_slv(x : int1736_t) return std_logic_vector;
function slv_to_int1736_t(x : std_logic_vector) return int1736_t;
subtype uint1737_t is unsigned(1736 downto 0);
constant uint1737_t_SLV_LEN : integer := 1737;
function uint1737_t_to_slv(x : uint1737_t) return std_logic_vector;
function slv_to_uint1737_t(x : std_logic_vector) return uint1737_t;
subtype int1737_t is signed(1736 downto 0);
constant int1737_t_SLV_LEN : integer := 1737;
function int1737_t_to_slv(x : int1737_t) return std_logic_vector;
function slv_to_int1737_t(x : std_logic_vector) return int1737_t;
subtype uint1738_t is unsigned(1737 downto 0);
constant uint1738_t_SLV_LEN : integer := 1738;
function uint1738_t_to_slv(x : uint1738_t) return std_logic_vector;
function slv_to_uint1738_t(x : std_logic_vector) return uint1738_t;
subtype int1738_t is signed(1737 downto 0);
constant int1738_t_SLV_LEN : integer := 1738;
function int1738_t_to_slv(x : int1738_t) return std_logic_vector;
function slv_to_int1738_t(x : std_logic_vector) return int1738_t;
subtype uint1739_t is unsigned(1738 downto 0);
constant uint1739_t_SLV_LEN : integer := 1739;
function uint1739_t_to_slv(x : uint1739_t) return std_logic_vector;
function slv_to_uint1739_t(x : std_logic_vector) return uint1739_t;
subtype int1739_t is signed(1738 downto 0);
constant int1739_t_SLV_LEN : integer := 1739;
function int1739_t_to_slv(x : int1739_t) return std_logic_vector;
function slv_to_int1739_t(x : std_logic_vector) return int1739_t;
subtype uint1740_t is unsigned(1739 downto 0);
constant uint1740_t_SLV_LEN : integer := 1740;
function uint1740_t_to_slv(x : uint1740_t) return std_logic_vector;
function slv_to_uint1740_t(x : std_logic_vector) return uint1740_t;
subtype int1740_t is signed(1739 downto 0);
constant int1740_t_SLV_LEN : integer := 1740;
function int1740_t_to_slv(x : int1740_t) return std_logic_vector;
function slv_to_int1740_t(x : std_logic_vector) return int1740_t;
subtype uint1741_t is unsigned(1740 downto 0);
constant uint1741_t_SLV_LEN : integer := 1741;
function uint1741_t_to_slv(x : uint1741_t) return std_logic_vector;
function slv_to_uint1741_t(x : std_logic_vector) return uint1741_t;
subtype int1741_t is signed(1740 downto 0);
constant int1741_t_SLV_LEN : integer := 1741;
function int1741_t_to_slv(x : int1741_t) return std_logic_vector;
function slv_to_int1741_t(x : std_logic_vector) return int1741_t;
subtype uint1742_t is unsigned(1741 downto 0);
constant uint1742_t_SLV_LEN : integer := 1742;
function uint1742_t_to_slv(x : uint1742_t) return std_logic_vector;
function slv_to_uint1742_t(x : std_logic_vector) return uint1742_t;
subtype int1742_t is signed(1741 downto 0);
constant int1742_t_SLV_LEN : integer := 1742;
function int1742_t_to_slv(x : int1742_t) return std_logic_vector;
function slv_to_int1742_t(x : std_logic_vector) return int1742_t;
subtype uint1743_t is unsigned(1742 downto 0);
constant uint1743_t_SLV_LEN : integer := 1743;
function uint1743_t_to_slv(x : uint1743_t) return std_logic_vector;
function slv_to_uint1743_t(x : std_logic_vector) return uint1743_t;
subtype int1743_t is signed(1742 downto 0);
constant int1743_t_SLV_LEN : integer := 1743;
function int1743_t_to_slv(x : int1743_t) return std_logic_vector;
function slv_to_int1743_t(x : std_logic_vector) return int1743_t;
subtype uint1744_t is unsigned(1743 downto 0);
constant uint1744_t_SLV_LEN : integer := 1744;
function uint1744_t_to_slv(x : uint1744_t) return std_logic_vector;
function slv_to_uint1744_t(x : std_logic_vector) return uint1744_t;
subtype int1744_t is signed(1743 downto 0);
constant int1744_t_SLV_LEN : integer := 1744;
function int1744_t_to_slv(x : int1744_t) return std_logic_vector;
function slv_to_int1744_t(x : std_logic_vector) return int1744_t;
subtype uint1745_t is unsigned(1744 downto 0);
constant uint1745_t_SLV_LEN : integer := 1745;
function uint1745_t_to_slv(x : uint1745_t) return std_logic_vector;
function slv_to_uint1745_t(x : std_logic_vector) return uint1745_t;
subtype int1745_t is signed(1744 downto 0);
constant int1745_t_SLV_LEN : integer := 1745;
function int1745_t_to_slv(x : int1745_t) return std_logic_vector;
function slv_to_int1745_t(x : std_logic_vector) return int1745_t;
subtype uint1746_t is unsigned(1745 downto 0);
constant uint1746_t_SLV_LEN : integer := 1746;
function uint1746_t_to_slv(x : uint1746_t) return std_logic_vector;
function slv_to_uint1746_t(x : std_logic_vector) return uint1746_t;
subtype int1746_t is signed(1745 downto 0);
constant int1746_t_SLV_LEN : integer := 1746;
function int1746_t_to_slv(x : int1746_t) return std_logic_vector;
function slv_to_int1746_t(x : std_logic_vector) return int1746_t;
subtype uint1747_t is unsigned(1746 downto 0);
constant uint1747_t_SLV_LEN : integer := 1747;
function uint1747_t_to_slv(x : uint1747_t) return std_logic_vector;
function slv_to_uint1747_t(x : std_logic_vector) return uint1747_t;
subtype int1747_t is signed(1746 downto 0);
constant int1747_t_SLV_LEN : integer := 1747;
function int1747_t_to_slv(x : int1747_t) return std_logic_vector;
function slv_to_int1747_t(x : std_logic_vector) return int1747_t;
subtype uint1748_t is unsigned(1747 downto 0);
constant uint1748_t_SLV_LEN : integer := 1748;
function uint1748_t_to_slv(x : uint1748_t) return std_logic_vector;
function slv_to_uint1748_t(x : std_logic_vector) return uint1748_t;
subtype int1748_t is signed(1747 downto 0);
constant int1748_t_SLV_LEN : integer := 1748;
function int1748_t_to_slv(x : int1748_t) return std_logic_vector;
function slv_to_int1748_t(x : std_logic_vector) return int1748_t;
subtype uint1749_t is unsigned(1748 downto 0);
constant uint1749_t_SLV_LEN : integer := 1749;
function uint1749_t_to_slv(x : uint1749_t) return std_logic_vector;
function slv_to_uint1749_t(x : std_logic_vector) return uint1749_t;
subtype int1749_t is signed(1748 downto 0);
constant int1749_t_SLV_LEN : integer := 1749;
function int1749_t_to_slv(x : int1749_t) return std_logic_vector;
function slv_to_int1749_t(x : std_logic_vector) return int1749_t;
subtype uint1750_t is unsigned(1749 downto 0);
constant uint1750_t_SLV_LEN : integer := 1750;
function uint1750_t_to_slv(x : uint1750_t) return std_logic_vector;
function slv_to_uint1750_t(x : std_logic_vector) return uint1750_t;
subtype int1750_t is signed(1749 downto 0);
constant int1750_t_SLV_LEN : integer := 1750;
function int1750_t_to_slv(x : int1750_t) return std_logic_vector;
function slv_to_int1750_t(x : std_logic_vector) return int1750_t;
subtype uint1751_t is unsigned(1750 downto 0);
constant uint1751_t_SLV_LEN : integer := 1751;
function uint1751_t_to_slv(x : uint1751_t) return std_logic_vector;
function slv_to_uint1751_t(x : std_logic_vector) return uint1751_t;
subtype int1751_t is signed(1750 downto 0);
constant int1751_t_SLV_LEN : integer := 1751;
function int1751_t_to_slv(x : int1751_t) return std_logic_vector;
function slv_to_int1751_t(x : std_logic_vector) return int1751_t;
subtype uint1752_t is unsigned(1751 downto 0);
constant uint1752_t_SLV_LEN : integer := 1752;
function uint1752_t_to_slv(x : uint1752_t) return std_logic_vector;
function slv_to_uint1752_t(x : std_logic_vector) return uint1752_t;
subtype int1752_t is signed(1751 downto 0);
constant int1752_t_SLV_LEN : integer := 1752;
function int1752_t_to_slv(x : int1752_t) return std_logic_vector;
function slv_to_int1752_t(x : std_logic_vector) return int1752_t;
subtype uint1753_t is unsigned(1752 downto 0);
constant uint1753_t_SLV_LEN : integer := 1753;
function uint1753_t_to_slv(x : uint1753_t) return std_logic_vector;
function slv_to_uint1753_t(x : std_logic_vector) return uint1753_t;
subtype int1753_t is signed(1752 downto 0);
constant int1753_t_SLV_LEN : integer := 1753;
function int1753_t_to_slv(x : int1753_t) return std_logic_vector;
function slv_to_int1753_t(x : std_logic_vector) return int1753_t;
subtype uint1754_t is unsigned(1753 downto 0);
constant uint1754_t_SLV_LEN : integer := 1754;
function uint1754_t_to_slv(x : uint1754_t) return std_logic_vector;
function slv_to_uint1754_t(x : std_logic_vector) return uint1754_t;
subtype int1754_t is signed(1753 downto 0);
constant int1754_t_SLV_LEN : integer := 1754;
function int1754_t_to_slv(x : int1754_t) return std_logic_vector;
function slv_to_int1754_t(x : std_logic_vector) return int1754_t;
subtype uint1755_t is unsigned(1754 downto 0);
constant uint1755_t_SLV_LEN : integer := 1755;
function uint1755_t_to_slv(x : uint1755_t) return std_logic_vector;
function slv_to_uint1755_t(x : std_logic_vector) return uint1755_t;
subtype int1755_t is signed(1754 downto 0);
constant int1755_t_SLV_LEN : integer := 1755;
function int1755_t_to_slv(x : int1755_t) return std_logic_vector;
function slv_to_int1755_t(x : std_logic_vector) return int1755_t;
subtype uint1756_t is unsigned(1755 downto 0);
constant uint1756_t_SLV_LEN : integer := 1756;
function uint1756_t_to_slv(x : uint1756_t) return std_logic_vector;
function slv_to_uint1756_t(x : std_logic_vector) return uint1756_t;
subtype int1756_t is signed(1755 downto 0);
constant int1756_t_SLV_LEN : integer := 1756;
function int1756_t_to_slv(x : int1756_t) return std_logic_vector;
function slv_to_int1756_t(x : std_logic_vector) return int1756_t;
subtype uint1757_t is unsigned(1756 downto 0);
constant uint1757_t_SLV_LEN : integer := 1757;
function uint1757_t_to_slv(x : uint1757_t) return std_logic_vector;
function slv_to_uint1757_t(x : std_logic_vector) return uint1757_t;
subtype int1757_t is signed(1756 downto 0);
constant int1757_t_SLV_LEN : integer := 1757;
function int1757_t_to_slv(x : int1757_t) return std_logic_vector;
function slv_to_int1757_t(x : std_logic_vector) return int1757_t;
subtype uint1758_t is unsigned(1757 downto 0);
constant uint1758_t_SLV_LEN : integer := 1758;
function uint1758_t_to_slv(x : uint1758_t) return std_logic_vector;
function slv_to_uint1758_t(x : std_logic_vector) return uint1758_t;
subtype int1758_t is signed(1757 downto 0);
constant int1758_t_SLV_LEN : integer := 1758;
function int1758_t_to_slv(x : int1758_t) return std_logic_vector;
function slv_to_int1758_t(x : std_logic_vector) return int1758_t;
subtype uint1759_t is unsigned(1758 downto 0);
constant uint1759_t_SLV_LEN : integer := 1759;
function uint1759_t_to_slv(x : uint1759_t) return std_logic_vector;
function slv_to_uint1759_t(x : std_logic_vector) return uint1759_t;
subtype int1759_t is signed(1758 downto 0);
constant int1759_t_SLV_LEN : integer := 1759;
function int1759_t_to_slv(x : int1759_t) return std_logic_vector;
function slv_to_int1759_t(x : std_logic_vector) return int1759_t;
subtype uint1760_t is unsigned(1759 downto 0);
constant uint1760_t_SLV_LEN : integer := 1760;
function uint1760_t_to_slv(x : uint1760_t) return std_logic_vector;
function slv_to_uint1760_t(x : std_logic_vector) return uint1760_t;
subtype int1760_t is signed(1759 downto 0);
constant int1760_t_SLV_LEN : integer := 1760;
function int1760_t_to_slv(x : int1760_t) return std_logic_vector;
function slv_to_int1760_t(x : std_logic_vector) return int1760_t;
subtype uint1761_t is unsigned(1760 downto 0);
constant uint1761_t_SLV_LEN : integer := 1761;
function uint1761_t_to_slv(x : uint1761_t) return std_logic_vector;
function slv_to_uint1761_t(x : std_logic_vector) return uint1761_t;
subtype int1761_t is signed(1760 downto 0);
constant int1761_t_SLV_LEN : integer := 1761;
function int1761_t_to_slv(x : int1761_t) return std_logic_vector;
function slv_to_int1761_t(x : std_logic_vector) return int1761_t;
subtype uint1762_t is unsigned(1761 downto 0);
constant uint1762_t_SLV_LEN : integer := 1762;
function uint1762_t_to_slv(x : uint1762_t) return std_logic_vector;
function slv_to_uint1762_t(x : std_logic_vector) return uint1762_t;
subtype int1762_t is signed(1761 downto 0);
constant int1762_t_SLV_LEN : integer := 1762;
function int1762_t_to_slv(x : int1762_t) return std_logic_vector;
function slv_to_int1762_t(x : std_logic_vector) return int1762_t;
subtype uint1763_t is unsigned(1762 downto 0);
constant uint1763_t_SLV_LEN : integer := 1763;
function uint1763_t_to_slv(x : uint1763_t) return std_logic_vector;
function slv_to_uint1763_t(x : std_logic_vector) return uint1763_t;
subtype int1763_t is signed(1762 downto 0);
constant int1763_t_SLV_LEN : integer := 1763;
function int1763_t_to_slv(x : int1763_t) return std_logic_vector;
function slv_to_int1763_t(x : std_logic_vector) return int1763_t;
subtype uint1764_t is unsigned(1763 downto 0);
constant uint1764_t_SLV_LEN : integer := 1764;
function uint1764_t_to_slv(x : uint1764_t) return std_logic_vector;
function slv_to_uint1764_t(x : std_logic_vector) return uint1764_t;
subtype int1764_t is signed(1763 downto 0);
constant int1764_t_SLV_LEN : integer := 1764;
function int1764_t_to_slv(x : int1764_t) return std_logic_vector;
function slv_to_int1764_t(x : std_logic_vector) return int1764_t;
subtype uint1765_t is unsigned(1764 downto 0);
constant uint1765_t_SLV_LEN : integer := 1765;
function uint1765_t_to_slv(x : uint1765_t) return std_logic_vector;
function slv_to_uint1765_t(x : std_logic_vector) return uint1765_t;
subtype int1765_t is signed(1764 downto 0);
constant int1765_t_SLV_LEN : integer := 1765;
function int1765_t_to_slv(x : int1765_t) return std_logic_vector;
function slv_to_int1765_t(x : std_logic_vector) return int1765_t;
subtype uint1766_t is unsigned(1765 downto 0);
constant uint1766_t_SLV_LEN : integer := 1766;
function uint1766_t_to_slv(x : uint1766_t) return std_logic_vector;
function slv_to_uint1766_t(x : std_logic_vector) return uint1766_t;
subtype int1766_t is signed(1765 downto 0);
constant int1766_t_SLV_LEN : integer := 1766;
function int1766_t_to_slv(x : int1766_t) return std_logic_vector;
function slv_to_int1766_t(x : std_logic_vector) return int1766_t;
subtype uint1767_t is unsigned(1766 downto 0);
constant uint1767_t_SLV_LEN : integer := 1767;
function uint1767_t_to_slv(x : uint1767_t) return std_logic_vector;
function slv_to_uint1767_t(x : std_logic_vector) return uint1767_t;
subtype int1767_t is signed(1766 downto 0);
constant int1767_t_SLV_LEN : integer := 1767;
function int1767_t_to_slv(x : int1767_t) return std_logic_vector;
function slv_to_int1767_t(x : std_logic_vector) return int1767_t;
subtype uint1768_t is unsigned(1767 downto 0);
constant uint1768_t_SLV_LEN : integer := 1768;
function uint1768_t_to_slv(x : uint1768_t) return std_logic_vector;
function slv_to_uint1768_t(x : std_logic_vector) return uint1768_t;
subtype int1768_t is signed(1767 downto 0);
constant int1768_t_SLV_LEN : integer := 1768;
function int1768_t_to_slv(x : int1768_t) return std_logic_vector;
function slv_to_int1768_t(x : std_logic_vector) return int1768_t;
subtype uint1769_t is unsigned(1768 downto 0);
constant uint1769_t_SLV_LEN : integer := 1769;
function uint1769_t_to_slv(x : uint1769_t) return std_logic_vector;
function slv_to_uint1769_t(x : std_logic_vector) return uint1769_t;
subtype int1769_t is signed(1768 downto 0);
constant int1769_t_SLV_LEN : integer := 1769;
function int1769_t_to_slv(x : int1769_t) return std_logic_vector;
function slv_to_int1769_t(x : std_logic_vector) return int1769_t;
subtype uint1770_t is unsigned(1769 downto 0);
constant uint1770_t_SLV_LEN : integer := 1770;
function uint1770_t_to_slv(x : uint1770_t) return std_logic_vector;
function slv_to_uint1770_t(x : std_logic_vector) return uint1770_t;
subtype int1770_t is signed(1769 downto 0);
constant int1770_t_SLV_LEN : integer := 1770;
function int1770_t_to_slv(x : int1770_t) return std_logic_vector;
function slv_to_int1770_t(x : std_logic_vector) return int1770_t;
subtype uint1771_t is unsigned(1770 downto 0);
constant uint1771_t_SLV_LEN : integer := 1771;
function uint1771_t_to_slv(x : uint1771_t) return std_logic_vector;
function slv_to_uint1771_t(x : std_logic_vector) return uint1771_t;
subtype int1771_t is signed(1770 downto 0);
constant int1771_t_SLV_LEN : integer := 1771;
function int1771_t_to_slv(x : int1771_t) return std_logic_vector;
function slv_to_int1771_t(x : std_logic_vector) return int1771_t;
subtype uint1772_t is unsigned(1771 downto 0);
constant uint1772_t_SLV_LEN : integer := 1772;
function uint1772_t_to_slv(x : uint1772_t) return std_logic_vector;
function slv_to_uint1772_t(x : std_logic_vector) return uint1772_t;
subtype int1772_t is signed(1771 downto 0);
constant int1772_t_SLV_LEN : integer := 1772;
function int1772_t_to_slv(x : int1772_t) return std_logic_vector;
function slv_to_int1772_t(x : std_logic_vector) return int1772_t;
subtype uint1773_t is unsigned(1772 downto 0);
constant uint1773_t_SLV_LEN : integer := 1773;
function uint1773_t_to_slv(x : uint1773_t) return std_logic_vector;
function slv_to_uint1773_t(x : std_logic_vector) return uint1773_t;
subtype int1773_t is signed(1772 downto 0);
constant int1773_t_SLV_LEN : integer := 1773;
function int1773_t_to_slv(x : int1773_t) return std_logic_vector;
function slv_to_int1773_t(x : std_logic_vector) return int1773_t;
subtype uint1774_t is unsigned(1773 downto 0);
constant uint1774_t_SLV_LEN : integer := 1774;
function uint1774_t_to_slv(x : uint1774_t) return std_logic_vector;
function slv_to_uint1774_t(x : std_logic_vector) return uint1774_t;
subtype int1774_t is signed(1773 downto 0);
constant int1774_t_SLV_LEN : integer := 1774;
function int1774_t_to_slv(x : int1774_t) return std_logic_vector;
function slv_to_int1774_t(x : std_logic_vector) return int1774_t;
subtype uint1775_t is unsigned(1774 downto 0);
constant uint1775_t_SLV_LEN : integer := 1775;
function uint1775_t_to_slv(x : uint1775_t) return std_logic_vector;
function slv_to_uint1775_t(x : std_logic_vector) return uint1775_t;
subtype int1775_t is signed(1774 downto 0);
constant int1775_t_SLV_LEN : integer := 1775;
function int1775_t_to_slv(x : int1775_t) return std_logic_vector;
function slv_to_int1775_t(x : std_logic_vector) return int1775_t;
subtype uint1776_t is unsigned(1775 downto 0);
constant uint1776_t_SLV_LEN : integer := 1776;
function uint1776_t_to_slv(x : uint1776_t) return std_logic_vector;
function slv_to_uint1776_t(x : std_logic_vector) return uint1776_t;
subtype int1776_t is signed(1775 downto 0);
constant int1776_t_SLV_LEN : integer := 1776;
function int1776_t_to_slv(x : int1776_t) return std_logic_vector;
function slv_to_int1776_t(x : std_logic_vector) return int1776_t;
subtype uint1777_t is unsigned(1776 downto 0);
constant uint1777_t_SLV_LEN : integer := 1777;
function uint1777_t_to_slv(x : uint1777_t) return std_logic_vector;
function slv_to_uint1777_t(x : std_logic_vector) return uint1777_t;
subtype int1777_t is signed(1776 downto 0);
constant int1777_t_SLV_LEN : integer := 1777;
function int1777_t_to_slv(x : int1777_t) return std_logic_vector;
function slv_to_int1777_t(x : std_logic_vector) return int1777_t;
subtype uint1778_t is unsigned(1777 downto 0);
constant uint1778_t_SLV_LEN : integer := 1778;
function uint1778_t_to_slv(x : uint1778_t) return std_logic_vector;
function slv_to_uint1778_t(x : std_logic_vector) return uint1778_t;
subtype int1778_t is signed(1777 downto 0);
constant int1778_t_SLV_LEN : integer := 1778;
function int1778_t_to_slv(x : int1778_t) return std_logic_vector;
function slv_to_int1778_t(x : std_logic_vector) return int1778_t;
subtype uint1779_t is unsigned(1778 downto 0);
constant uint1779_t_SLV_LEN : integer := 1779;
function uint1779_t_to_slv(x : uint1779_t) return std_logic_vector;
function slv_to_uint1779_t(x : std_logic_vector) return uint1779_t;
subtype int1779_t is signed(1778 downto 0);
constant int1779_t_SLV_LEN : integer := 1779;
function int1779_t_to_slv(x : int1779_t) return std_logic_vector;
function slv_to_int1779_t(x : std_logic_vector) return int1779_t;
subtype uint1780_t is unsigned(1779 downto 0);
constant uint1780_t_SLV_LEN : integer := 1780;
function uint1780_t_to_slv(x : uint1780_t) return std_logic_vector;
function slv_to_uint1780_t(x : std_logic_vector) return uint1780_t;
subtype int1780_t is signed(1779 downto 0);
constant int1780_t_SLV_LEN : integer := 1780;
function int1780_t_to_slv(x : int1780_t) return std_logic_vector;
function slv_to_int1780_t(x : std_logic_vector) return int1780_t;
subtype uint1781_t is unsigned(1780 downto 0);
constant uint1781_t_SLV_LEN : integer := 1781;
function uint1781_t_to_slv(x : uint1781_t) return std_logic_vector;
function slv_to_uint1781_t(x : std_logic_vector) return uint1781_t;
subtype int1781_t is signed(1780 downto 0);
constant int1781_t_SLV_LEN : integer := 1781;
function int1781_t_to_slv(x : int1781_t) return std_logic_vector;
function slv_to_int1781_t(x : std_logic_vector) return int1781_t;
subtype uint1782_t is unsigned(1781 downto 0);
constant uint1782_t_SLV_LEN : integer := 1782;
function uint1782_t_to_slv(x : uint1782_t) return std_logic_vector;
function slv_to_uint1782_t(x : std_logic_vector) return uint1782_t;
subtype int1782_t is signed(1781 downto 0);
constant int1782_t_SLV_LEN : integer := 1782;
function int1782_t_to_slv(x : int1782_t) return std_logic_vector;
function slv_to_int1782_t(x : std_logic_vector) return int1782_t;
subtype uint1783_t is unsigned(1782 downto 0);
constant uint1783_t_SLV_LEN : integer := 1783;
function uint1783_t_to_slv(x : uint1783_t) return std_logic_vector;
function slv_to_uint1783_t(x : std_logic_vector) return uint1783_t;
subtype int1783_t is signed(1782 downto 0);
constant int1783_t_SLV_LEN : integer := 1783;
function int1783_t_to_slv(x : int1783_t) return std_logic_vector;
function slv_to_int1783_t(x : std_logic_vector) return int1783_t;
subtype uint1784_t is unsigned(1783 downto 0);
constant uint1784_t_SLV_LEN : integer := 1784;
function uint1784_t_to_slv(x : uint1784_t) return std_logic_vector;
function slv_to_uint1784_t(x : std_logic_vector) return uint1784_t;
subtype int1784_t is signed(1783 downto 0);
constant int1784_t_SLV_LEN : integer := 1784;
function int1784_t_to_slv(x : int1784_t) return std_logic_vector;
function slv_to_int1784_t(x : std_logic_vector) return int1784_t;
subtype uint1785_t is unsigned(1784 downto 0);
constant uint1785_t_SLV_LEN : integer := 1785;
function uint1785_t_to_slv(x : uint1785_t) return std_logic_vector;
function slv_to_uint1785_t(x : std_logic_vector) return uint1785_t;
subtype int1785_t is signed(1784 downto 0);
constant int1785_t_SLV_LEN : integer := 1785;
function int1785_t_to_slv(x : int1785_t) return std_logic_vector;
function slv_to_int1785_t(x : std_logic_vector) return int1785_t;
subtype uint1786_t is unsigned(1785 downto 0);
constant uint1786_t_SLV_LEN : integer := 1786;
function uint1786_t_to_slv(x : uint1786_t) return std_logic_vector;
function slv_to_uint1786_t(x : std_logic_vector) return uint1786_t;
subtype int1786_t is signed(1785 downto 0);
constant int1786_t_SLV_LEN : integer := 1786;
function int1786_t_to_slv(x : int1786_t) return std_logic_vector;
function slv_to_int1786_t(x : std_logic_vector) return int1786_t;
subtype uint1787_t is unsigned(1786 downto 0);
constant uint1787_t_SLV_LEN : integer := 1787;
function uint1787_t_to_slv(x : uint1787_t) return std_logic_vector;
function slv_to_uint1787_t(x : std_logic_vector) return uint1787_t;
subtype int1787_t is signed(1786 downto 0);
constant int1787_t_SLV_LEN : integer := 1787;
function int1787_t_to_slv(x : int1787_t) return std_logic_vector;
function slv_to_int1787_t(x : std_logic_vector) return int1787_t;
subtype uint1788_t is unsigned(1787 downto 0);
constant uint1788_t_SLV_LEN : integer := 1788;
function uint1788_t_to_slv(x : uint1788_t) return std_logic_vector;
function slv_to_uint1788_t(x : std_logic_vector) return uint1788_t;
subtype int1788_t is signed(1787 downto 0);
constant int1788_t_SLV_LEN : integer := 1788;
function int1788_t_to_slv(x : int1788_t) return std_logic_vector;
function slv_to_int1788_t(x : std_logic_vector) return int1788_t;
subtype uint1789_t is unsigned(1788 downto 0);
constant uint1789_t_SLV_LEN : integer := 1789;
function uint1789_t_to_slv(x : uint1789_t) return std_logic_vector;
function slv_to_uint1789_t(x : std_logic_vector) return uint1789_t;
subtype int1789_t is signed(1788 downto 0);
constant int1789_t_SLV_LEN : integer := 1789;
function int1789_t_to_slv(x : int1789_t) return std_logic_vector;
function slv_to_int1789_t(x : std_logic_vector) return int1789_t;
subtype uint1790_t is unsigned(1789 downto 0);
constant uint1790_t_SLV_LEN : integer := 1790;
function uint1790_t_to_slv(x : uint1790_t) return std_logic_vector;
function slv_to_uint1790_t(x : std_logic_vector) return uint1790_t;
subtype int1790_t is signed(1789 downto 0);
constant int1790_t_SLV_LEN : integer := 1790;
function int1790_t_to_slv(x : int1790_t) return std_logic_vector;
function slv_to_int1790_t(x : std_logic_vector) return int1790_t;
subtype uint1791_t is unsigned(1790 downto 0);
constant uint1791_t_SLV_LEN : integer := 1791;
function uint1791_t_to_slv(x : uint1791_t) return std_logic_vector;
function slv_to_uint1791_t(x : std_logic_vector) return uint1791_t;
subtype int1791_t is signed(1790 downto 0);
constant int1791_t_SLV_LEN : integer := 1791;
function int1791_t_to_slv(x : int1791_t) return std_logic_vector;
function slv_to_int1791_t(x : std_logic_vector) return int1791_t;
subtype uint1792_t is unsigned(1791 downto 0);
constant uint1792_t_SLV_LEN : integer := 1792;
function uint1792_t_to_slv(x : uint1792_t) return std_logic_vector;
function slv_to_uint1792_t(x : std_logic_vector) return uint1792_t;
subtype int1792_t is signed(1791 downto 0);
constant int1792_t_SLV_LEN : integer := 1792;
function int1792_t_to_slv(x : int1792_t) return std_logic_vector;
function slv_to_int1792_t(x : std_logic_vector) return int1792_t;
subtype uint1793_t is unsigned(1792 downto 0);
constant uint1793_t_SLV_LEN : integer := 1793;
function uint1793_t_to_slv(x : uint1793_t) return std_logic_vector;
function slv_to_uint1793_t(x : std_logic_vector) return uint1793_t;
subtype int1793_t is signed(1792 downto 0);
constant int1793_t_SLV_LEN : integer := 1793;
function int1793_t_to_slv(x : int1793_t) return std_logic_vector;
function slv_to_int1793_t(x : std_logic_vector) return int1793_t;
subtype uint1794_t is unsigned(1793 downto 0);
constant uint1794_t_SLV_LEN : integer := 1794;
function uint1794_t_to_slv(x : uint1794_t) return std_logic_vector;
function slv_to_uint1794_t(x : std_logic_vector) return uint1794_t;
subtype int1794_t is signed(1793 downto 0);
constant int1794_t_SLV_LEN : integer := 1794;
function int1794_t_to_slv(x : int1794_t) return std_logic_vector;
function slv_to_int1794_t(x : std_logic_vector) return int1794_t;
subtype uint1795_t is unsigned(1794 downto 0);
constant uint1795_t_SLV_LEN : integer := 1795;
function uint1795_t_to_slv(x : uint1795_t) return std_logic_vector;
function slv_to_uint1795_t(x : std_logic_vector) return uint1795_t;
subtype int1795_t is signed(1794 downto 0);
constant int1795_t_SLV_LEN : integer := 1795;
function int1795_t_to_slv(x : int1795_t) return std_logic_vector;
function slv_to_int1795_t(x : std_logic_vector) return int1795_t;
subtype uint1796_t is unsigned(1795 downto 0);
constant uint1796_t_SLV_LEN : integer := 1796;
function uint1796_t_to_slv(x : uint1796_t) return std_logic_vector;
function slv_to_uint1796_t(x : std_logic_vector) return uint1796_t;
subtype int1796_t is signed(1795 downto 0);
constant int1796_t_SLV_LEN : integer := 1796;
function int1796_t_to_slv(x : int1796_t) return std_logic_vector;
function slv_to_int1796_t(x : std_logic_vector) return int1796_t;
subtype uint1797_t is unsigned(1796 downto 0);
constant uint1797_t_SLV_LEN : integer := 1797;
function uint1797_t_to_slv(x : uint1797_t) return std_logic_vector;
function slv_to_uint1797_t(x : std_logic_vector) return uint1797_t;
subtype int1797_t is signed(1796 downto 0);
constant int1797_t_SLV_LEN : integer := 1797;
function int1797_t_to_slv(x : int1797_t) return std_logic_vector;
function slv_to_int1797_t(x : std_logic_vector) return int1797_t;
subtype uint1798_t is unsigned(1797 downto 0);
constant uint1798_t_SLV_LEN : integer := 1798;
function uint1798_t_to_slv(x : uint1798_t) return std_logic_vector;
function slv_to_uint1798_t(x : std_logic_vector) return uint1798_t;
subtype int1798_t is signed(1797 downto 0);
constant int1798_t_SLV_LEN : integer := 1798;
function int1798_t_to_slv(x : int1798_t) return std_logic_vector;
function slv_to_int1798_t(x : std_logic_vector) return int1798_t;
subtype uint1799_t is unsigned(1798 downto 0);
constant uint1799_t_SLV_LEN : integer := 1799;
function uint1799_t_to_slv(x : uint1799_t) return std_logic_vector;
function slv_to_uint1799_t(x : std_logic_vector) return uint1799_t;
subtype int1799_t is signed(1798 downto 0);
constant int1799_t_SLV_LEN : integer := 1799;
function int1799_t_to_slv(x : int1799_t) return std_logic_vector;
function slv_to_int1799_t(x : std_logic_vector) return int1799_t;
subtype uint1800_t is unsigned(1799 downto 0);
constant uint1800_t_SLV_LEN : integer := 1800;
function uint1800_t_to_slv(x : uint1800_t) return std_logic_vector;
function slv_to_uint1800_t(x : std_logic_vector) return uint1800_t;
subtype int1800_t is signed(1799 downto 0);
constant int1800_t_SLV_LEN : integer := 1800;
function int1800_t_to_slv(x : int1800_t) return std_logic_vector;
function slv_to_int1800_t(x : std_logic_vector) return int1800_t;
subtype uint1801_t is unsigned(1800 downto 0);
constant uint1801_t_SLV_LEN : integer := 1801;
function uint1801_t_to_slv(x : uint1801_t) return std_logic_vector;
function slv_to_uint1801_t(x : std_logic_vector) return uint1801_t;
subtype int1801_t is signed(1800 downto 0);
constant int1801_t_SLV_LEN : integer := 1801;
function int1801_t_to_slv(x : int1801_t) return std_logic_vector;
function slv_to_int1801_t(x : std_logic_vector) return int1801_t;
subtype uint1802_t is unsigned(1801 downto 0);
constant uint1802_t_SLV_LEN : integer := 1802;
function uint1802_t_to_slv(x : uint1802_t) return std_logic_vector;
function slv_to_uint1802_t(x : std_logic_vector) return uint1802_t;
subtype int1802_t is signed(1801 downto 0);
constant int1802_t_SLV_LEN : integer := 1802;
function int1802_t_to_slv(x : int1802_t) return std_logic_vector;
function slv_to_int1802_t(x : std_logic_vector) return int1802_t;
subtype uint1803_t is unsigned(1802 downto 0);
constant uint1803_t_SLV_LEN : integer := 1803;
function uint1803_t_to_slv(x : uint1803_t) return std_logic_vector;
function slv_to_uint1803_t(x : std_logic_vector) return uint1803_t;
subtype int1803_t is signed(1802 downto 0);
constant int1803_t_SLV_LEN : integer := 1803;
function int1803_t_to_slv(x : int1803_t) return std_logic_vector;
function slv_to_int1803_t(x : std_logic_vector) return int1803_t;
subtype uint1804_t is unsigned(1803 downto 0);
constant uint1804_t_SLV_LEN : integer := 1804;
function uint1804_t_to_slv(x : uint1804_t) return std_logic_vector;
function slv_to_uint1804_t(x : std_logic_vector) return uint1804_t;
subtype int1804_t is signed(1803 downto 0);
constant int1804_t_SLV_LEN : integer := 1804;
function int1804_t_to_slv(x : int1804_t) return std_logic_vector;
function slv_to_int1804_t(x : std_logic_vector) return int1804_t;
subtype uint1805_t is unsigned(1804 downto 0);
constant uint1805_t_SLV_LEN : integer := 1805;
function uint1805_t_to_slv(x : uint1805_t) return std_logic_vector;
function slv_to_uint1805_t(x : std_logic_vector) return uint1805_t;
subtype int1805_t is signed(1804 downto 0);
constant int1805_t_SLV_LEN : integer := 1805;
function int1805_t_to_slv(x : int1805_t) return std_logic_vector;
function slv_to_int1805_t(x : std_logic_vector) return int1805_t;
subtype uint1806_t is unsigned(1805 downto 0);
constant uint1806_t_SLV_LEN : integer := 1806;
function uint1806_t_to_slv(x : uint1806_t) return std_logic_vector;
function slv_to_uint1806_t(x : std_logic_vector) return uint1806_t;
subtype int1806_t is signed(1805 downto 0);
constant int1806_t_SLV_LEN : integer := 1806;
function int1806_t_to_slv(x : int1806_t) return std_logic_vector;
function slv_to_int1806_t(x : std_logic_vector) return int1806_t;
subtype uint1807_t is unsigned(1806 downto 0);
constant uint1807_t_SLV_LEN : integer := 1807;
function uint1807_t_to_slv(x : uint1807_t) return std_logic_vector;
function slv_to_uint1807_t(x : std_logic_vector) return uint1807_t;
subtype int1807_t is signed(1806 downto 0);
constant int1807_t_SLV_LEN : integer := 1807;
function int1807_t_to_slv(x : int1807_t) return std_logic_vector;
function slv_to_int1807_t(x : std_logic_vector) return int1807_t;
subtype uint1808_t is unsigned(1807 downto 0);
constant uint1808_t_SLV_LEN : integer := 1808;
function uint1808_t_to_slv(x : uint1808_t) return std_logic_vector;
function slv_to_uint1808_t(x : std_logic_vector) return uint1808_t;
subtype int1808_t is signed(1807 downto 0);
constant int1808_t_SLV_LEN : integer := 1808;
function int1808_t_to_slv(x : int1808_t) return std_logic_vector;
function slv_to_int1808_t(x : std_logic_vector) return int1808_t;
subtype uint1809_t is unsigned(1808 downto 0);
constant uint1809_t_SLV_LEN : integer := 1809;
function uint1809_t_to_slv(x : uint1809_t) return std_logic_vector;
function slv_to_uint1809_t(x : std_logic_vector) return uint1809_t;
subtype int1809_t is signed(1808 downto 0);
constant int1809_t_SLV_LEN : integer := 1809;
function int1809_t_to_slv(x : int1809_t) return std_logic_vector;
function slv_to_int1809_t(x : std_logic_vector) return int1809_t;
subtype uint1810_t is unsigned(1809 downto 0);
constant uint1810_t_SLV_LEN : integer := 1810;
function uint1810_t_to_slv(x : uint1810_t) return std_logic_vector;
function slv_to_uint1810_t(x : std_logic_vector) return uint1810_t;
subtype int1810_t is signed(1809 downto 0);
constant int1810_t_SLV_LEN : integer := 1810;
function int1810_t_to_slv(x : int1810_t) return std_logic_vector;
function slv_to_int1810_t(x : std_logic_vector) return int1810_t;
subtype uint1811_t is unsigned(1810 downto 0);
constant uint1811_t_SLV_LEN : integer := 1811;
function uint1811_t_to_slv(x : uint1811_t) return std_logic_vector;
function slv_to_uint1811_t(x : std_logic_vector) return uint1811_t;
subtype int1811_t is signed(1810 downto 0);
constant int1811_t_SLV_LEN : integer := 1811;
function int1811_t_to_slv(x : int1811_t) return std_logic_vector;
function slv_to_int1811_t(x : std_logic_vector) return int1811_t;
subtype uint1812_t is unsigned(1811 downto 0);
constant uint1812_t_SLV_LEN : integer := 1812;
function uint1812_t_to_slv(x : uint1812_t) return std_logic_vector;
function slv_to_uint1812_t(x : std_logic_vector) return uint1812_t;
subtype int1812_t is signed(1811 downto 0);
constant int1812_t_SLV_LEN : integer := 1812;
function int1812_t_to_slv(x : int1812_t) return std_logic_vector;
function slv_to_int1812_t(x : std_logic_vector) return int1812_t;
subtype uint1813_t is unsigned(1812 downto 0);
constant uint1813_t_SLV_LEN : integer := 1813;
function uint1813_t_to_slv(x : uint1813_t) return std_logic_vector;
function slv_to_uint1813_t(x : std_logic_vector) return uint1813_t;
subtype int1813_t is signed(1812 downto 0);
constant int1813_t_SLV_LEN : integer := 1813;
function int1813_t_to_slv(x : int1813_t) return std_logic_vector;
function slv_to_int1813_t(x : std_logic_vector) return int1813_t;
subtype uint1814_t is unsigned(1813 downto 0);
constant uint1814_t_SLV_LEN : integer := 1814;
function uint1814_t_to_slv(x : uint1814_t) return std_logic_vector;
function slv_to_uint1814_t(x : std_logic_vector) return uint1814_t;
subtype int1814_t is signed(1813 downto 0);
constant int1814_t_SLV_LEN : integer := 1814;
function int1814_t_to_slv(x : int1814_t) return std_logic_vector;
function slv_to_int1814_t(x : std_logic_vector) return int1814_t;
subtype uint1815_t is unsigned(1814 downto 0);
constant uint1815_t_SLV_LEN : integer := 1815;
function uint1815_t_to_slv(x : uint1815_t) return std_logic_vector;
function slv_to_uint1815_t(x : std_logic_vector) return uint1815_t;
subtype int1815_t is signed(1814 downto 0);
constant int1815_t_SLV_LEN : integer := 1815;
function int1815_t_to_slv(x : int1815_t) return std_logic_vector;
function slv_to_int1815_t(x : std_logic_vector) return int1815_t;
subtype uint1816_t is unsigned(1815 downto 0);
constant uint1816_t_SLV_LEN : integer := 1816;
function uint1816_t_to_slv(x : uint1816_t) return std_logic_vector;
function slv_to_uint1816_t(x : std_logic_vector) return uint1816_t;
subtype int1816_t is signed(1815 downto 0);
constant int1816_t_SLV_LEN : integer := 1816;
function int1816_t_to_slv(x : int1816_t) return std_logic_vector;
function slv_to_int1816_t(x : std_logic_vector) return int1816_t;
subtype uint1817_t is unsigned(1816 downto 0);
constant uint1817_t_SLV_LEN : integer := 1817;
function uint1817_t_to_slv(x : uint1817_t) return std_logic_vector;
function slv_to_uint1817_t(x : std_logic_vector) return uint1817_t;
subtype int1817_t is signed(1816 downto 0);
constant int1817_t_SLV_LEN : integer := 1817;
function int1817_t_to_slv(x : int1817_t) return std_logic_vector;
function slv_to_int1817_t(x : std_logic_vector) return int1817_t;
subtype uint1818_t is unsigned(1817 downto 0);
constant uint1818_t_SLV_LEN : integer := 1818;
function uint1818_t_to_slv(x : uint1818_t) return std_logic_vector;
function slv_to_uint1818_t(x : std_logic_vector) return uint1818_t;
subtype int1818_t is signed(1817 downto 0);
constant int1818_t_SLV_LEN : integer := 1818;
function int1818_t_to_slv(x : int1818_t) return std_logic_vector;
function slv_to_int1818_t(x : std_logic_vector) return int1818_t;
subtype uint1819_t is unsigned(1818 downto 0);
constant uint1819_t_SLV_LEN : integer := 1819;
function uint1819_t_to_slv(x : uint1819_t) return std_logic_vector;
function slv_to_uint1819_t(x : std_logic_vector) return uint1819_t;
subtype int1819_t is signed(1818 downto 0);
constant int1819_t_SLV_LEN : integer := 1819;
function int1819_t_to_slv(x : int1819_t) return std_logic_vector;
function slv_to_int1819_t(x : std_logic_vector) return int1819_t;
subtype uint1820_t is unsigned(1819 downto 0);
constant uint1820_t_SLV_LEN : integer := 1820;
function uint1820_t_to_slv(x : uint1820_t) return std_logic_vector;
function slv_to_uint1820_t(x : std_logic_vector) return uint1820_t;
subtype int1820_t is signed(1819 downto 0);
constant int1820_t_SLV_LEN : integer := 1820;
function int1820_t_to_slv(x : int1820_t) return std_logic_vector;
function slv_to_int1820_t(x : std_logic_vector) return int1820_t;
subtype uint1821_t is unsigned(1820 downto 0);
constant uint1821_t_SLV_LEN : integer := 1821;
function uint1821_t_to_slv(x : uint1821_t) return std_logic_vector;
function slv_to_uint1821_t(x : std_logic_vector) return uint1821_t;
subtype int1821_t is signed(1820 downto 0);
constant int1821_t_SLV_LEN : integer := 1821;
function int1821_t_to_slv(x : int1821_t) return std_logic_vector;
function slv_to_int1821_t(x : std_logic_vector) return int1821_t;
subtype uint1822_t is unsigned(1821 downto 0);
constant uint1822_t_SLV_LEN : integer := 1822;
function uint1822_t_to_slv(x : uint1822_t) return std_logic_vector;
function slv_to_uint1822_t(x : std_logic_vector) return uint1822_t;
subtype int1822_t is signed(1821 downto 0);
constant int1822_t_SLV_LEN : integer := 1822;
function int1822_t_to_slv(x : int1822_t) return std_logic_vector;
function slv_to_int1822_t(x : std_logic_vector) return int1822_t;
subtype uint1823_t is unsigned(1822 downto 0);
constant uint1823_t_SLV_LEN : integer := 1823;
function uint1823_t_to_slv(x : uint1823_t) return std_logic_vector;
function slv_to_uint1823_t(x : std_logic_vector) return uint1823_t;
subtype int1823_t is signed(1822 downto 0);
constant int1823_t_SLV_LEN : integer := 1823;
function int1823_t_to_slv(x : int1823_t) return std_logic_vector;
function slv_to_int1823_t(x : std_logic_vector) return int1823_t;
subtype uint1824_t is unsigned(1823 downto 0);
constant uint1824_t_SLV_LEN : integer := 1824;
function uint1824_t_to_slv(x : uint1824_t) return std_logic_vector;
function slv_to_uint1824_t(x : std_logic_vector) return uint1824_t;
subtype int1824_t is signed(1823 downto 0);
constant int1824_t_SLV_LEN : integer := 1824;
function int1824_t_to_slv(x : int1824_t) return std_logic_vector;
function slv_to_int1824_t(x : std_logic_vector) return int1824_t;
subtype uint1825_t is unsigned(1824 downto 0);
constant uint1825_t_SLV_LEN : integer := 1825;
function uint1825_t_to_slv(x : uint1825_t) return std_logic_vector;
function slv_to_uint1825_t(x : std_logic_vector) return uint1825_t;
subtype int1825_t is signed(1824 downto 0);
constant int1825_t_SLV_LEN : integer := 1825;
function int1825_t_to_slv(x : int1825_t) return std_logic_vector;
function slv_to_int1825_t(x : std_logic_vector) return int1825_t;
subtype uint1826_t is unsigned(1825 downto 0);
constant uint1826_t_SLV_LEN : integer := 1826;
function uint1826_t_to_slv(x : uint1826_t) return std_logic_vector;
function slv_to_uint1826_t(x : std_logic_vector) return uint1826_t;
subtype int1826_t is signed(1825 downto 0);
constant int1826_t_SLV_LEN : integer := 1826;
function int1826_t_to_slv(x : int1826_t) return std_logic_vector;
function slv_to_int1826_t(x : std_logic_vector) return int1826_t;
subtype uint1827_t is unsigned(1826 downto 0);
constant uint1827_t_SLV_LEN : integer := 1827;
function uint1827_t_to_slv(x : uint1827_t) return std_logic_vector;
function slv_to_uint1827_t(x : std_logic_vector) return uint1827_t;
subtype int1827_t is signed(1826 downto 0);
constant int1827_t_SLV_LEN : integer := 1827;
function int1827_t_to_slv(x : int1827_t) return std_logic_vector;
function slv_to_int1827_t(x : std_logic_vector) return int1827_t;
subtype uint1828_t is unsigned(1827 downto 0);
constant uint1828_t_SLV_LEN : integer := 1828;
function uint1828_t_to_slv(x : uint1828_t) return std_logic_vector;
function slv_to_uint1828_t(x : std_logic_vector) return uint1828_t;
subtype int1828_t is signed(1827 downto 0);
constant int1828_t_SLV_LEN : integer := 1828;
function int1828_t_to_slv(x : int1828_t) return std_logic_vector;
function slv_to_int1828_t(x : std_logic_vector) return int1828_t;
subtype uint1829_t is unsigned(1828 downto 0);
constant uint1829_t_SLV_LEN : integer := 1829;
function uint1829_t_to_slv(x : uint1829_t) return std_logic_vector;
function slv_to_uint1829_t(x : std_logic_vector) return uint1829_t;
subtype int1829_t is signed(1828 downto 0);
constant int1829_t_SLV_LEN : integer := 1829;
function int1829_t_to_slv(x : int1829_t) return std_logic_vector;
function slv_to_int1829_t(x : std_logic_vector) return int1829_t;
subtype uint1830_t is unsigned(1829 downto 0);
constant uint1830_t_SLV_LEN : integer := 1830;
function uint1830_t_to_slv(x : uint1830_t) return std_logic_vector;
function slv_to_uint1830_t(x : std_logic_vector) return uint1830_t;
subtype int1830_t is signed(1829 downto 0);
constant int1830_t_SLV_LEN : integer := 1830;
function int1830_t_to_slv(x : int1830_t) return std_logic_vector;
function slv_to_int1830_t(x : std_logic_vector) return int1830_t;
subtype uint1831_t is unsigned(1830 downto 0);
constant uint1831_t_SLV_LEN : integer := 1831;
function uint1831_t_to_slv(x : uint1831_t) return std_logic_vector;
function slv_to_uint1831_t(x : std_logic_vector) return uint1831_t;
subtype int1831_t is signed(1830 downto 0);
constant int1831_t_SLV_LEN : integer := 1831;
function int1831_t_to_slv(x : int1831_t) return std_logic_vector;
function slv_to_int1831_t(x : std_logic_vector) return int1831_t;
subtype uint1832_t is unsigned(1831 downto 0);
constant uint1832_t_SLV_LEN : integer := 1832;
function uint1832_t_to_slv(x : uint1832_t) return std_logic_vector;
function slv_to_uint1832_t(x : std_logic_vector) return uint1832_t;
subtype int1832_t is signed(1831 downto 0);
constant int1832_t_SLV_LEN : integer := 1832;
function int1832_t_to_slv(x : int1832_t) return std_logic_vector;
function slv_to_int1832_t(x : std_logic_vector) return int1832_t;
subtype uint1833_t is unsigned(1832 downto 0);
constant uint1833_t_SLV_LEN : integer := 1833;
function uint1833_t_to_slv(x : uint1833_t) return std_logic_vector;
function slv_to_uint1833_t(x : std_logic_vector) return uint1833_t;
subtype int1833_t is signed(1832 downto 0);
constant int1833_t_SLV_LEN : integer := 1833;
function int1833_t_to_slv(x : int1833_t) return std_logic_vector;
function slv_to_int1833_t(x : std_logic_vector) return int1833_t;
subtype uint1834_t is unsigned(1833 downto 0);
constant uint1834_t_SLV_LEN : integer := 1834;
function uint1834_t_to_slv(x : uint1834_t) return std_logic_vector;
function slv_to_uint1834_t(x : std_logic_vector) return uint1834_t;
subtype int1834_t is signed(1833 downto 0);
constant int1834_t_SLV_LEN : integer := 1834;
function int1834_t_to_slv(x : int1834_t) return std_logic_vector;
function slv_to_int1834_t(x : std_logic_vector) return int1834_t;
subtype uint1835_t is unsigned(1834 downto 0);
constant uint1835_t_SLV_LEN : integer := 1835;
function uint1835_t_to_slv(x : uint1835_t) return std_logic_vector;
function slv_to_uint1835_t(x : std_logic_vector) return uint1835_t;
subtype int1835_t is signed(1834 downto 0);
constant int1835_t_SLV_LEN : integer := 1835;
function int1835_t_to_slv(x : int1835_t) return std_logic_vector;
function slv_to_int1835_t(x : std_logic_vector) return int1835_t;
subtype uint1836_t is unsigned(1835 downto 0);
constant uint1836_t_SLV_LEN : integer := 1836;
function uint1836_t_to_slv(x : uint1836_t) return std_logic_vector;
function slv_to_uint1836_t(x : std_logic_vector) return uint1836_t;
subtype int1836_t is signed(1835 downto 0);
constant int1836_t_SLV_LEN : integer := 1836;
function int1836_t_to_slv(x : int1836_t) return std_logic_vector;
function slv_to_int1836_t(x : std_logic_vector) return int1836_t;
subtype uint1837_t is unsigned(1836 downto 0);
constant uint1837_t_SLV_LEN : integer := 1837;
function uint1837_t_to_slv(x : uint1837_t) return std_logic_vector;
function slv_to_uint1837_t(x : std_logic_vector) return uint1837_t;
subtype int1837_t is signed(1836 downto 0);
constant int1837_t_SLV_LEN : integer := 1837;
function int1837_t_to_slv(x : int1837_t) return std_logic_vector;
function slv_to_int1837_t(x : std_logic_vector) return int1837_t;
subtype uint1838_t is unsigned(1837 downto 0);
constant uint1838_t_SLV_LEN : integer := 1838;
function uint1838_t_to_slv(x : uint1838_t) return std_logic_vector;
function slv_to_uint1838_t(x : std_logic_vector) return uint1838_t;
subtype int1838_t is signed(1837 downto 0);
constant int1838_t_SLV_LEN : integer := 1838;
function int1838_t_to_slv(x : int1838_t) return std_logic_vector;
function slv_to_int1838_t(x : std_logic_vector) return int1838_t;
subtype uint1839_t is unsigned(1838 downto 0);
constant uint1839_t_SLV_LEN : integer := 1839;
function uint1839_t_to_slv(x : uint1839_t) return std_logic_vector;
function slv_to_uint1839_t(x : std_logic_vector) return uint1839_t;
subtype int1839_t is signed(1838 downto 0);
constant int1839_t_SLV_LEN : integer := 1839;
function int1839_t_to_slv(x : int1839_t) return std_logic_vector;
function slv_to_int1839_t(x : std_logic_vector) return int1839_t;
subtype uint1840_t is unsigned(1839 downto 0);
constant uint1840_t_SLV_LEN : integer := 1840;
function uint1840_t_to_slv(x : uint1840_t) return std_logic_vector;
function slv_to_uint1840_t(x : std_logic_vector) return uint1840_t;
subtype int1840_t is signed(1839 downto 0);
constant int1840_t_SLV_LEN : integer := 1840;
function int1840_t_to_slv(x : int1840_t) return std_logic_vector;
function slv_to_int1840_t(x : std_logic_vector) return int1840_t;
subtype uint1841_t is unsigned(1840 downto 0);
constant uint1841_t_SLV_LEN : integer := 1841;
function uint1841_t_to_slv(x : uint1841_t) return std_logic_vector;
function slv_to_uint1841_t(x : std_logic_vector) return uint1841_t;
subtype int1841_t is signed(1840 downto 0);
constant int1841_t_SLV_LEN : integer := 1841;
function int1841_t_to_slv(x : int1841_t) return std_logic_vector;
function slv_to_int1841_t(x : std_logic_vector) return int1841_t;
subtype uint1842_t is unsigned(1841 downto 0);
constant uint1842_t_SLV_LEN : integer := 1842;
function uint1842_t_to_slv(x : uint1842_t) return std_logic_vector;
function slv_to_uint1842_t(x : std_logic_vector) return uint1842_t;
subtype int1842_t is signed(1841 downto 0);
constant int1842_t_SLV_LEN : integer := 1842;
function int1842_t_to_slv(x : int1842_t) return std_logic_vector;
function slv_to_int1842_t(x : std_logic_vector) return int1842_t;
subtype uint1843_t is unsigned(1842 downto 0);
constant uint1843_t_SLV_LEN : integer := 1843;
function uint1843_t_to_slv(x : uint1843_t) return std_logic_vector;
function slv_to_uint1843_t(x : std_logic_vector) return uint1843_t;
subtype int1843_t is signed(1842 downto 0);
constant int1843_t_SLV_LEN : integer := 1843;
function int1843_t_to_slv(x : int1843_t) return std_logic_vector;
function slv_to_int1843_t(x : std_logic_vector) return int1843_t;
subtype uint1844_t is unsigned(1843 downto 0);
constant uint1844_t_SLV_LEN : integer := 1844;
function uint1844_t_to_slv(x : uint1844_t) return std_logic_vector;
function slv_to_uint1844_t(x : std_logic_vector) return uint1844_t;
subtype int1844_t is signed(1843 downto 0);
constant int1844_t_SLV_LEN : integer := 1844;
function int1844_t_to_slv(x : int1844_t) return std_logic_vector;
function slv_to_int1844_t(x : std_logic_vector) return int1844_t;
subtype uint1845_t is unsigned(1844 downto 0);
constant uint1845_t_SLV_LEN : integer := 1845;
function uint1845_t_to_slv(x : uint1845_t) return std_logic_vector;
function slv_to_uint1845_t(x : std_logic_vector) return uint1845_t;
subtype int1845_t is signed(1844 downto 0);
constant int1845_t_SLV_LEN : integer := 1845;
function int1845_t_to_slv(x : int1845_t) return std_logic_vector;
function slv_to_int1845_t(x : std_logic_vector) return int1845_t;
subtype uint1846_t is unsigned(1845 downto 0);
constant uint1846_t_SLV_LEN : integer := 1846;
function uint1846_t_to_slv(x : uint1846_t) return std_logic_vector;
function slv_to_uint1846_t(x : std_logic_vector) return uint1846_t;
subtype int1846_t is signed(1845 downto 0);
constant int1846_t_SLV_LEN : integer := 1846;
function int1846_t_to_slv(x : int1846_t) return std_logic_vector;
function slv_to_int1846_t(x : std_logic_vector) return int1846_t;
subtype uint1847_t is unsigned(1846 downto 0);
constant uint1847_t_SLV_LEN : integer := 1847;
function uint1847_t_to_slv(x : uint1847_t) return std_logic_vector;
function slv_to_uint1847_t(x : std_logic_vector) return uint1847_t;
subtype int1847_t is signed(1846 downto 0);
constant int1847_t_SLV_LEN : integer := 1847;
function int1847_t_to_slv(x : int1847_t) return std_logic_vector;
function slv_to_int1847_t(x : std_logic_vector) return int1847_t;
subtype uint1848_t is unsigned(1847 downto 0);
constant uint1848_t_SLV_LEN : integer := 1848;
function uint1848_t_to_slv(x : uint1848_t) return std_logic_vector;
function slv_to_uint1848_t(x : std_logic_vector) return uint1848_t;
subtype int1848_t is signed(1847 downto 0);
constant int1848_t_SLV_LEN : integer := 1848;
function int1848_t_to_slv(x : int1848_t) return std_logic_vector;
function slv_to_int1848_t(x : std_logic_vector) return int1848_t;
subtype uint1849_t is unsigned(1848 downto 0);
constant uint1849_t_SLV_LEN : integer := 1849;
function uint1849_t_to_slv(x : uint1849_t) return std_logic_vector;
function slv_to_uint1849_t(x : std_logic_vector) return uint1849_t;
subtype int1849_t is signed(1848 downto 0);
constant int1849_t_SLV_LEN : integer := 1849;
function int1849_t_to_slv(x : int1849_t) return std_logic_vector;
function slv_to_int1849_t(x : std_logic_vector) return int1849_t;
subtype uint1850_t is unsigned(1849 downto 0);
constant uint1850_t_SLV_LEN : integer := 1850;
function uint1850_t_to_slv(x : uint1850_t) return std_logic_vector;
function slv_to_uint1850_t(x : std_logic_vector) return uint1850_t;
subtype int1850_t is signed(1849 downto 0);
constant int1850_t_SLV_LEN : integer := 1850;
function int1850_t_to_slv(x : int1850_t) return std_logic_vector;
function slv_to_int1850_t(x : std_logic_vector) return int1850_t;
subtype uint1851_t is unsigned(1850 downto 0);
constant uint1851_t_SLV_LEN : integer := 1851;
function uint1851_t_to_slv(x : uint1851_t) return std_logic_vector;
function slv_to_uint1851_t(x : std_logic_vector) return uint1851_t;
subtype int1851_t is signed(1850 downto 0);
constant int1851_t_SLV_LEN : integer := 1851;
function int1851_t_to_slv(x : int1851_t) return std_logic_vector;
function slv_to_int1851_t(x : std_logic_vector) return int1851_t;
subtype uint1852_t is unsigned(1851 downto 0);
constant uint1852_t_SLV_LEN : integer := 1852;
function uint1852_t_to_slv(x : uint1852_t) return std_logic_vector;
function slv_to_uint1852_t(x : std_logic_vector) return uint1852_t;
subtype int1852_t is signed(1851 downto 0);
constant int1852_t_SLV_LEN : integer := 1852;
function int1852_t_to_slv(x : int1852_t) return std_logic_vector;
function slv_to_int1852_t(x : std_logic_vector) return int1852_t;
subtype uint1853_t is unsigned(1852 downto 0);
constant uint1853_t_SLV_LEN : integer := 1853;
function uint1853_t_to_slv(x : uint1853_t) return std_logic_vector;
function slv_to_uint1853_t(x : std_logic_vector) return uint1853_t;
subtype int1853_t is signed(1852 downto 0);
constant int1853_t_SLV_LEN : integer := 1853;
function int1853_t_to_slv(x : int1853_t) return std_logic_vector;
function slv_to_int1853_t(x : std_logic_vector) return int1853_t;
subtype uint1854_t is unsigned(1853 downto 0);
constant uint1854_t_SLV_LEN : integer := 1854;
function uint1854_t_to_slv(x : uint1854_t) return std_logic_vector;
function slv_to_uint1854_t(x : std_logic_vector) return uint1854_t;
subtype int1854_t is signed(1853 downto 0);
constant int1854_t_SLV_LEN : integer := 1854;
function int1854_t_to_slv(x : int1854_t) return std_logic_vector;
function slv_to_int1854_t(x : std_logic_vector) return int1854_t;
subtype uint1855_t is unsigned(1854 downto 0);
constant uint1855_t_SLV_LEN : integer := 1855;
function uint1855_t_to_slv(x : uint1855_t) return std_logic_vector;
function slv_to_uint1855_t(x : std_logic_vector) return uint1855_t;
subtype int1855_t is signed(1854 downto 0);
constant int1855_t_SLV_LEN : integer := 1855;
function int1855_t_to_slv(x : int1855_t) return std_logic_vector;
function slv_to_int1855_t(x : std_logic_vector) return int1855_t;
subtype uint1856_t is unsigned(1855 downto 0);
constant uint1856_t_SLV_LEN : integer := 1856;
function uint1856_t_to_slv(x : uint1856_t) return std_logic_vector;
function slv_to_uint1856_t(x : std_logic_vector) return uint1856_t;
subtype int1856_t is signed(1855 downto 0);
constant int1856_t_SLV_LEN : integer := 1856;
function int1856_t_to_slv(x : int1856_t) return std_logic_vector;
function slv_to_int1856_t(x : std_logic_vector) return int1856_t;
subtype uint1857_t is unsigned(1856 downto 0);
constant uint1857_t_SLV_LEN : integer := 1857;
function uint1857_t_to_slv(x : uint1857_t) return std_logic_vector;
function slv_to_uint1857_t(x : std_logic_vector) return uint1857_t;
subtype int1857_t is signed(1856 downto 0);
constant int1857_t_SLV_LEN : integer := 1857;
function int1857_t_to_slv(x : int1857_t) return std_logic_vector;
function slv_to_int1857_t(x : std_logic_vector) return int1857_t;
subtype uint1858_t is unsigned(1857 downto 0);
constant uint1858_t_SLV_LEN : integer := 1858;
function uint1858_t_to_slv(x : uint1858_t) return std_logic_vector;
function slv_to_uint1858_t(x : std_logic_vector) return uint1858_t;
subtype int1858_t is signed(1857 downto 0);
constant int1858_t_SLV_LEN : integer := 1858;
function int1858_t_to_slv(x : int1858_t) return std_logic_vector;
function slv_to_int1858_t(x : std_logic_vector) return int1858_t;
subtype uint1859_t is unsigned(1858 downto 0);
constant uint1859_t_SLV_LEN : integer := 1859;
function uint1859_t_to_slv(x : uint1859_t) return std_logic_vector;
function slv_to_uint1859_t(x : std_logic_vector) return uint1859_t;
subtype int1859_t is signed(1858 downto 0);
constant int1859_t_SLV_LEN : integer := 1859;
function int1859_t_to_slv(x : int1859_t) return std_logic_vector;
function slv_to_int1859_t(x : std_logic_vector) return int1859_t;
subtype uint1860_t is unsigned(1859 downto 0);
constant uint1860_t_SLV_LEN : integer := 1860;
function uint1860_t_to_slv(x : uint1860_t) return std_logic_vector;
function slv_to_uint1860_t(x : std_logic_vector) return uint1860_t;
subtype int1860_t is signed(1859 downto 0);
constant int1860_t_SLV_LEN : integer := 1860;
function int1860_t_to_slv(x : int1860_t) return std_logic_vector;
function slv_to_int1860_t(x : std_logic_vector) return int1860_t;
subtype uint1861_t is unsigned(1860 downto 0);
constant uint1861_t_SLV_LEN : integer := 1861;
function uint1861_t_to_slv(x : uint1861_t) return std_logic_vector;
function slv_to_uint1861_t(x : std_logic_vector) return uint1861_t;
subtype int1861_t is signed(1860 downto 0);
constant int1861_t_SLV_LEN : integer := 1861;
function int1861_t_to_slv(x : int1861_t) return std_logic_vector;
function slv_to_int1861_t(x : std_logic_vector) return int1861_t;
subtype uint1862_t is unsigned(1861 downto 0);
constant uint1862_t_SLV_LEN : integer := 1862;
function uint1862_t_to_slv(x : uint1862_t) return std_logic_vector;
function slv_to_uint1862_t(x : std_logic_vector) return uint1862_t;
subtype int1862_t is signed(1861 downto 0);
constant int1862_t_SLV_LEN : integer := 1862;
function int1862_t_to_slv(x : int1862_t) return std_logic_vector;
function slv_to_int1862_t(x : std_logic_vector) return int1862_t;
subtype uint1863_t is unsigned(1862 downto 0);
constant uint1863_t_SLV_LEN : integer := 1863;
function uint1863_t_to_slv(x : uint1863_t) return std_logic_vector;
function slv_to_uint1863_t(x : std_logic_vector) return uint1863_t;
subtype int1863_t is signed(1862 downto 0);
constant int1863_t_SLV_LEN : integer := 1863;
function int1863_t_to_slv(x : int1863_t) return std_logic_vector;
function slv_to_int1863_t(x : std_logic_vector) return int1863_t;
subtype uint1864_t is unsigned(1863 downto 0);
constant uint1864_t_SLV_LEN : integer := 1864;
function uint1864_t_to_slv(x : uint1864_t) return std_logic_vector;
function slv_to_uint1864_t(x : std_logic_vector) return uint1864_t;
subtype int1864_t is signed(1863 downto 0);
constant int1864_t_SLV_LEN : integer := 1864;
function int1864_t_to_slv(x : int1864_t) return std_logic_vector;
function slv_to_int1864_t(x : std_logic_vector) return int1864_t;
subtype uint1865_t is unsigned(1864 downto 0);
constant uint1865_t_SLV_LEN : integer := 1865;
function uint1865_t_to_slv(x : uint1865_t) return std_logic_vector;
function slv_to_uint1865_t(x : std_logic_vector) return uint1865_t;
subtype int1865_t is signed(1864 downto 0);
constant int1865_t_SLV_LEN : integer := 1865;
function int1865_t_to_slv(x : int1865_t) return std_logic_vector;
function slv_to_int1865_t(x : std_logic_vector) return int1865_t;
subtype uint1866_t is unsigned(1865 downto 0);
constant uint1866_t_SLV_LEN : integer := 1866;
function uint1866_t_to_slv(x : uint1866_t) return std_logic_vector;
function slv_to_uint1866_t(x : std_logic_vector) return uint1866_t;
subtype int1866_t is signed(1865 downto 0);
constant int1866_t_SLV_LEN : integer := 1866;
function int1866_t_to_slv(x : int1866_t) return std_logic_vector;
function slv_to_int1866_t(x : std_logic_vector) return int1866_t;
subtype uint1867_t is unsigned(1866 downto 0);
constant uint1867_t_SLV_LEN : integer := 1867;
function uint1867_t_to_slv(x : uint1867_t) return std_logic_vector;
function slv_to_uint1867_t(x : std_logic_vector) return uint1867_t;
subtype int1867_t is signed(1866 downto 0);
constant int1867_t_SLV_LEN : integer := 1867;
function int1867_t_to_slv(x : int1867_t) return std_logic_vector;
function slv_to_int1867_t(x : std_logic_vector) return int1867_t;
subtype uint1868_t is unsigned(1867 downto 0);
constant uint1868_t_SLV_LEN : integer := 1868;
function uint1868_t_to_slv(x : uint1868_t) return std_logic_vector;
function slv_to_uint1868_t(x : std_logic_vector) return uint1868_t;
subtype int1868_t is signed(1867 downto 0);
constant int1868_t_SLV_LEN : integer := 1868;
function int1868_t_to_slv(x : int1868_t) return std_logic_vector;
function slv_to_int1868_t(x : std_logic_vector) return int1868_t;
subtype uint1869_t is unsigned(1868 downto 0);
constant uint1869_t_SLV_LEN : integer := 1869;
function uint1869_t_to_slv(x : uint1869_t) return std_logic_vector;
function slv_to_uint1869_t(x : std_logic_vector) return uint1869_t;
subtype int1869_t is signed(1868 downto 0);
constant int1869_t_SLV_LEN : integer := 1869;
function int1869_t_to_slv(x : int1869_t) return std_logic_vector;
function slv_to_int1869_t(x : std_logic_vector) return int1869_t;
subtype uint1870_t is unsigned(1869 downto 0);
constant uint1870_t_SLV_LEN : integer := 1870;
function uint1870_t_to_slv(x : uint1870_t) return std_logic_vector;
function slv_to_uint1870_t(x : std_logic_vector) return uint1870_t;
subtype int1870_t is signed(1869 downto 0);
constant int1870_t_SLV_LEN : integer := 1870;
function int1870_t_to_slv(x : int1870_t) return std_logic_vector;
function slv_to_int1870_t(x : std_logic_vector) return int1870_t;
subtype uint1871_t is unsigned(1870 downto 0);
constant uint1871_t_SLV_LEN : integer := 1871;
function uint1871_t_to_slv(x : uint1871_t) return std_logic_vector;
function slv_to_uint1871_t(x : std_logic_vector) return uint1871_t;
subtype int1871_t is signed(1870 downto 0);
constant int1871_t_SLV_LEN : integer := 1871;
function int1871_t_to_slv(x : int1871_t) return std_logic_vector;
function slv_to_int1871_t(x : std_logic_vector) return int1871_t;
subtype uint1872_t is unsigned(1871 downto 0);
constant uint1872_t_SLV_LEN : integer := 1872;
function uint1872_t_to_slv(x : uint1872_t) return std_logic_vector;
function slv_to_uint1872_t(x : std_logic_vector) return uint1872_t;
subtype int1872_t is signed(1871 downto 0);
constant int1872_t_SLV_LEN : integer := 1872;
function int1872_t_to_slv(x : int1872_t) return std_logic_vector;
function slv_to_int1872_t(x : std_logic_vector) return int1872_t;
subtype uint1873_t is unsigned(1872 downto 0);
constant uint1873_t_SLV_LEN : integer := 1873;
function uint1873_t_to_slv(x : uint1873_t) return std_logic_vector;
function slv_to_uint1873_t(x : std_logic_vector) return uint1873_t;
subtype int1873_t is signed(1872 downto 0);
constant int1873_t_SLV_LEN : integer := 1873;
function int1873_t_to_slv(x : int1873_t) return std_logic_vector;
function slv_to_int1873_t(x : std_logic_vector) return int1873_t;
subtype uint1874_t is unsigned(1873 downto 0);
constant uint1874_t_SLV_LEN : integer := 1874;
function uint1874_t_to_slv(x : uint1874_t) return std_logic_vector;
function slv_to_uint1874_t(x : std_logic_vector) return uint1874_t;
subtype int1874_t is signed(1873 downto 0);
constant int1874_t_SLV_LEN : integer := 1874;
function int1874_t_to_slv(x : int1874_t) return std_logic_vector;
function slv_to_int1874_t(x : std_logic_vector) return int1874_t;
subtype uint1875_t is unsigned(1874 downto 0);
constant uint1875_t_SLV_LEN : integer := 1875;
function uint1875_t_to_slv(x : uint1875_t) return std_logic_vector;
function slv_to_uint1875_t(x : std_logic_vector) return uint1875_t;
subtype int1875_t is signed(1874 downto 0);
constant int1875_t_SLV_LEN : integer := 1875;
function int1875_t_to_slv(x : int1875_t) return std_logic_vector;
function slv_to_int1875_t(x : std_logic_vector) return int1875_t;
subtype uint1876_t is unsigned(1875 downto 0);
constant uint1876_t_SLV_LEN : integer := 1876;
function uint1876_t_to_slv(x : uint1876_t) return std_logic_vector;
function slv_to_uint1876_t(x : std_logic_vector) return uint1876_t;
subtype int1876_t is signed(1875 downto 0);
constant int1876_t_SLV_LEN : integer := 1876;
function int1876_t_to_slv(x : int1876_t) return std_logic_vector;
function slv_to_int1876_t(x : std_logic_vector) return int1876_t;
subtype uint1877_t is unsigned(1876 downto 0);
constant uint1877_t_SLV_LEN : integer := 1877;
function uint1877_t_to_slv(x : uint1877_t) return std_logic_vector;
function slv_to_uint1877_t(x : std_logic_vector) return uint1877_t;
subtype int1877_t is signed(1876 downto 0);
constant int1877_t_SLV_LEN : integer := 1877;
function int1877_t_to_slv(x : int1877_t) return std_logic_vector;
function slv_to_int1877_t(x : std_logic_vector) return int1877_t;
subtype uint1878_t is unsigned(1877 downto 0);
constant uint1878_t_SLV_LEN : integer := 1878;
function uint1878_t_to_slv(x : uint1878_t) return std_logic_vector;
function slv_to_uint1878_t(x : std_logic_vector) return uint1878_t;
subtype int1878_t is signed(1877 downto 0);
constant int1878_t_SLV_LEN : integer := 1878;
function int1878_t_to_slv(x : int1878_t) return std_logic_vector;
function slv_to_int1878_t(x : std_logic_vector) return int1878_t;
subtype uint1879_t is unsigned(1878 downto 0);
constant uint1879_t_SLV_LEN : integer := 1879;
function uint1879_t_to_slv(x : uint1879_t) return std_logic_vector;
function slv_to_uint1879_t(x : std_logic_vector) return uint1879_t;
subtype int1879_t is signed(1878 downto 0);
constant int1879_t_SLV_LEN : integer := 1879;
function int1879_t_to_slv(x : int1879_t) return std_logic_vector;
function slv_to_int1879_t(x : std_logic_vector) return int1879_t;
subtype uint1880_t is unsigned(1879 downto 0);
constant uint1880_t_SLV_LEN : integer := 1880;
function uint1880_t_to_slv(x : uint1880_t) return std_logic_vector;
function slv_to_uint1880_t(x : std_logic_vector) return uint1880_t;
subtype int1880_t is signed(1879 downto 0);
constant int1880_t_SLV_LEN : integer := 1880;
function int1880_t_to_slv(x : int1880_t) return std_logic_vector;
function slv_to_int1880_t(x : std_logic_vector) return int1880_t;
subtype uint1881_t is unsigned(1880 downto 0);
constant uint1881_t_SLV_LEN : integer := 1881;
function uint1881_t_to_slv(x : uint1881_t) return std_logic_vector;
function slv_to_uint1881_t(x : std_logic_vector) return uint1881_t;
subtype int1881_t is signed(1880 downto 0);
constant int1881_t_SLV_LEN : integer := 1881;
function int1881_t_to_slv(x : int1881_t) return std_logic_vector;
function slv_to_int1881_t(x : std_logic_vector) return int1881_t;
subtype uint1882_t is unsigned(1881 downto 0);
constant uint1882_t_SLV_LEN : integer := 1882;
function uint1882_t_to_slv(x : uint1882_t) return std_logic_vector;
function slv_to_uint1882_t(x : std_logic_vector) return uint1882_t;
subtype int1882_t is signed(1881 downto 0);
constant int1882_t_SLV_LEN : integer := 1882;
function int1882_t_to_slv(x : int1882_t) return std_logic_vector;
function slv_to_int1882_t(x : std_logic_vector) return int1882_t;
subtype uint1883_t is unsigned(1882 downto 0);
constant uint1883_t_SLV_LEN : integer := 1883;
function uint1883_t_to_slv(x : uint1883_t) return std_logic_vector;
function slv_to_uint1883_t(x : std_logic_vector) return uint1883_t;
subtype int1883_t is signed(1882 downto 0);
constant int1883_t_SLV_LEN : integer := 1883;
function int1883_t_to_slv(x : int1883_t) return std_logic_vector;
function slv_to_int1883_t(x : std_logic_vector) return int1883_t;
subtype uint1884_t is unsigned(1883 downto 0);
constant uint1884_t_SLV_LEN : integer := 1884;
function uint1884_t_to_slv(x : uint1884_t) return std_logic_vector;
function slv_to_uint1884_t(x : std_logic_vector) return uint1884_t;
subtype int1884_t is signed(1883 downto 0);
constant int1884_t_SLV_LEN : integer := 1884;
function int1884_t_to_slv(x : int1884_t) return std_logic_vector;
function slv_to_int1884_t(x : std_logic_vector) return int1884_t;
subtype uint1885_t is unsigned(1884 downto 0);
constant uint1885_t_SLV_LEN : integer := 1885;
function uint1885_t_to_slv(x : uint1885_t) return std_logic_vector;
function slv_to_uint1885_t(x : std_logic_vector) return uint1885_t;
subtype int1885_t is signed(1884 downto 0);
constant int1885_t_SLV_LEN : integer := 1885;
function int1885_t_to_slv(x : int1885_t) return std_logic_vector;
function slv_to_int1885_t(x : std_logic_vector) return int1885_t;
subtype uint1886_t is unsigned(1885 downto 0);
constant uint1886_t_SLV_LEN : integer := 1886;
function uint1886_t_to_slv(x : uint1886_t) return std_logic_vector;
function slv_to_uint1886_t(x : std_logic_vector) return uint1886_t;
subtype int1886_t is signed(1885 downto 0);
constant int1886_t_SLV_LEN : integer := 1886;
function int1886_t_to_slv(x : int1886_t) return std_logic_vector;
function slv_to_int1886_t(x : std_logic_vector) return int1886_t;
subtype uint1887_t is unsigned(1886 downto 0);
constant uint1887_t_SLV_LEN : integer := 1887;
function uint1887_t_to_slv(x : uint1887_t) return std_logic_vector;
function slv_to_uint1887_t(x : std_logic_vector) return uint1887_t;
subtype int1887_t is signed(1886 downto 0);
constant int1887_t_SLV_LEN : integer := 1887;
function int1887_t_to_slv(x : int1887_t) return std_logic_vector;
function slv_to_int1887_t(x : std_logic_vector) return int1887_t;
subtype uint1888_t is unsigned(1887 downto 0);
constant uint1888_t_SLV_LEN : integer := 1888;
function uint1888_t_to_slv(x : uint1888_t) return std_logic_vector;
function slv_to_uint1888_t(x : std_logic_vector) return uint1888_t;
subtype int1888_t is signed(1887 downto 0);
constant int1888_t_SLV_LEN : integer := 1888;
function int1888_t_to_slv(x : int1888_t) return std_logic_vector;
function slv_to_int1888_t(x : std_logic_vector) return int1888_t;
subtype uint1889_t is unsigned(1888 downto 0);
constant uint1889_t_SLV_LEN : integer := 1889;
function uint1889_t_to_slv(x : uint1889_t) return std_logic_vector;
function slv_to_uint1889_t(x : std_logic_vector) return uint1889_t;
subtype int1889_t is signed(1888 downto 0);
constant int1889_t_SLV_LEN : integer := 1889;
function int1889_t_to_slv(x : int1889_t) return std_logic_vector;
function slv_to_int1889_t(x : std_logic_vector) return int1889_t;
subtype uint1890_t is unsigned(1889 downto 0);
constant uint1890_t_SLV_LEN : integer := 1890;
function uint1890_t_to_slv(x : uint1890_t) return std_logic_vector;
function slv_to_uint1890_t(x : std_logic_vector) return uint1890_t;
subtype int1890_t is signed(1889 downto 0);
constant int1890_t_SLV_LEN : integer := 1890;
function int1890_t_to_slv(x : int1890_t) return std_logic_vector;
function slv_to_int1890_t(x : std_logic_vector) return int1890_t;
subtype uint1891_t is unsigned(1890 downto 0);
constant uint1891_t_SLV_LEN : integer := 1891;
function uint1891_t_to_slv(x : uint1891_t) return std_logic_vector;
function slv_to_uint1891_t(x : std_logic_vector) return uint1891_t;
subtype int1891_t is signed(1890 downto 0);
constant int1891_t_SLV_LEN : integer := 1891;
function int1891_t_to_slv(x : int1891_t) return std_logic_vector;
function slv_to_int1891_t(x : std_logic_vector) return int1891_t;
subtype uint1892_t is unsigned(1891 downto 0);
constant uint1892_t_SLV_LEN : integer := 1892;
function uint1892_t_to_slv(x : uint1892_t) return std_logic_vector;
function slv_to_uint1892_t(x : std_logic_vector) return uint1892_t;
subtype int1892_t is signed(1891 downto 0);
constant int1892_t_SLV_LEN : integer := 1892;
function int1892_t_to_slv(x : int1892_t) return std_logic_vector;
function slv_to_int1892_t(x : std_logic_vector) return int1892_t;
subtype uint1893_t is unsigned(1892 downto 0);
constant uint1893_t_SLV_LEN : integer := 1893;
function uint1893_t_to_slv(x : uint1893_t) return std_logic_vector;
function slv_to_uint1893_t(x : std_logic_vector) return uint1893_t;
subtype int1893_t is signed(1892 downto 0);
constant int1893_t_SLV_LEN : integer := 1893;
function int1893_t_to_slv(x : int1893_t) return std_logic_vector;
function slv_to_int1893_t(x : std_logic_vector) return int1893_t;
subtype uint1894_t is unsigned(1893 downto 0);
constant uint1894_t_SLV_LEN : integer := 1894;
function uint1894_t_to_slv(x : uint1894_t) return std_logic_vector;
function slv_to_uint1894_t(x : std_logic_vector) return uint1894_t;
subtype int1894_t is signed(1893 downto 0);
constant int1894_t_SLV_LEN : integer := 1894;
function int1894_t_to_slv(x : int1894_t) return std_logic_vector;
function slv_to_int1894_t(x : std_logic_vector) return int1894_t;
subtype uint1895_t is unsigned(1894 downto 0);
constant uint1895_t_SLV_LEN : integer := 1895;
function uint1895_t_to_slv(x : uint1895_t) return std_logic_vector;
function slv_to_uint1895_t(x : std_logic_vector) return uint1895_t;
subtype int1895_t is signed(1894 downto 0);
constant int1895_t_SLV_LEN : integer := 1895;
function int1895_t_to_slv(x : int1895_t) return std_logic_vector;
function slv_to_int1895_t(x : std_logic_vector) return int1895_t;
subtype uint1896_t is unsigned(1895 downto 0);
constant uint1896_t_SLV_LEN : integer := 1896;
function uint1896_t_to_slv(x : uint1896_t) return std_logic_vector;
function slv_to_uint1896_t(x : std_logic_vector) return uint1896_t;
subtype int1896_t is signed(1895 downto 0);
constant int1896_t_SLV_LEN : integer := 1896;
function int1896_t_to_slv(x : int1896_t) return std_logic_vector;
function slv_to_int1896_t(x : std_logic_vector) return int1896_t;
subtype uint1897_t is unsigned(1896 downto 0);
constant uint1897_t_SLV_LEN : integer := 1897;
function uint1897_t_to_slv(x : uint1897_t) return std_logic_vector;
function slv_to_uint1897_t(x : std_logic_vector) return uint1897_t;
subtype int1897_t is signed(1896 downto 0);
constant int1897_t_SLV_LEN : integer := 1897;
function int1897_t_to_slv(x : int1897_t) return std_logic_vector;
function slv_to_int1897_t(x : std_logic_vector) return int1897_t;
subtype uint1898_t is unsigned(1897 downto 0);
constant uint1898_t_SLV_LEN : integer := 1898;
function uint1898_t_to_slv(x : uint1898_t) return std_logic_vector;
function slv_to_uint1898_t(x : std_logic_vector) return uint1898_t;
subtype int1898_t is signed(1897 downto 0);
constant int1898_t_SLV_LEN : integer := 1898;
function int1898_t_to_slv(x : int1898_t) return std_logic_vector;
function slv_to_int1898_t(x : std_logic_vector) return int1898_t;
subtype uint1899_t is unsigned(1898 downto 0);
constant uint1899_t_SLV_LEN : integer := 1899;
function uint1899_t_to_slv(x : uint1899_t) return std_logic_vector;
function slv_to_uint1899_t(x : std_logic_vector) return uint1899_t;
subtype int1899_t is signed(1898 downto 0);
constant int1899_t_SLV_LEN : integer := 1899;
function int1899_t_to_slv(x : int1899_t) return std_logic_vector;
function slv_to_int1899_t(x : std_logic_vector) return int1899_t;
subtype uint1900_t is unsigned(1899 downto 0);
constant uint1900_t_SLV_LEN : integer := 1900;
function uint1900_t_to_slv(x : uint1900_t) return std_logic_vector;
function slv_to_uint1900_t(x : std_logic_vector) return uint1900_t;
subtype int1900_t is signed(1899 downto 0);
constant int1900_t_SLV_LEN : integer := 1900;
function int1900_t_to_slv(x : int1900_t) return std_logic_vector;
function slv_to_int1900_t(x : std_logic_vector) return int1900_t;
subtype uint1901_t is unsigned(1900 downto 0);
constant uint1901_t_SLV_LEN : integer := 1901;
function uint1901_t_to_slv(x : uint1901_t) return std_logic_vector;
function slv_to_uint1901_t(x : std_logic_vector) return uint1901_t;
subtype int1901_t is signed(1900 downto 0);
constant int1901_t_SLV_LEN : integer := 1901;
function int1901_t_to_slv(x : int1901_t) return std_logic_vector;
function slv_to_int1901_t(x : std_logic_vector) return int1901_t;
subtype uint1902_t is unsigned(1901 downto 0);
constant uint1902_t_SLV_LEN : integer := 1902;
function uint1902_t_to_slv(x : uint1902_t) return std_logic_vector;
function slv_to_uint1902_t(x : std_logic_vector) return uint1902_t;
subtype int1902_t is signed(1901 downto 0);
constant int1902_t_SLV_LEN : integer := 1902;
function int1902_t_to_slv(x : int1902_t) return std_logic_vector;
function slv_to_int1902_t(x : std_logic_vector) return int1902_t;
subtype uint1903_t is unsigned(1902 downto 0);
constant uint1903_t_SLV_LEN : integer := 1903;
function uint1903_t_to_slv(x : uint1903_t) return std_logic_vector;
function slv_to_uint1903_t(x : std_logic_vector) return uint1903_t;
subtype int1903_t is signed(1902 downto 0);
constant int1903_t_SLV_LEN : integer := 1903;
function int1903_t_to_slv(x : int1903_t) return std_logic_vector;
function slv_to_int1903_t(x : std_logic_vector) return int1903_t;
subtype uint1904_t is unsigned(1903 downto 0);
constant uint1904_t_SLV_LEN : integer := 1904;
function uint1904_t_to_slv(x : uint1904_t) return std_logic_vector;
function slv_to_uint1904_t(x : std_logic_vector) return uint1904_t;
subtype int1904_t is signed(1903 downto 0);
constant int1904_t_SLV_LEN : integer := 1904;
function int1904_t_to_slv(x : int1904_t) return std_logic_vector;
function slv_to_int1904_t(x : std_logic_vector) return int1904_t;
subtype uint1905_t is unsigned(1904 downto 0);
constant uint1905_t_SLV_LEN : integer := 1905;
function uint1905_t_to_slv(x : uint1905_t) return std_logic_vector;
function slv_to_uint1905_t(x : std_logic_vector) return uint1905_t;
subtype int1905_t is signed(1904 downto 0);
constant int1905_t_SLV_LEN : integer := 1905;
function int1905_t_to_slv(x : int1905_t) return std_logic_vector;
function slv_to_int1905_t(x : std_logic_vector) return int1905_t;
subtype uint1906_t is unsigned(1905 downto 0);
constant uint1906_t_SLV_LEN : integer := 1906;
function uint1906_t_to_slv(x : uint1906_t) return std_logic_vector;
function slv_to_uint1906_t(x : std_logic_vector) return uint1906_t;
subtype int1906_t is signed(1905 downto 0);
constant int1906_t_SLV_LEN : integer := 1906;
function int1906_t_to_slv(x : int1906_t) return std_logic_vector;
function slv_to_int1906_t(x : std_logic_vector) return int1906_t;
subtype uint1907_t is unsigned(1906 downto 0);
constant uint1907_t_SLV_LEN : integer := 1907;
function uint1907_t_to_slv(x : uint1907_t) return std_logic_vector;
function slv_to_uint1907_t(x : std_logic_vector) return uint1907_t;
subtype int1907_t is signed(1906 downto 0);
constant int1907_t_SLV_LEN : integer := 1907;
function int1907_t_to_slv(x : int1907_t) return std_logic_vector;
function slv_to_int1907_t(x : std_logic_vector) return int1907_t;
subtype uint1908_t is unsigned(1907 downto 0);
constant uint1908_t_SLV_LEN : integer := 1908;
function uint1908_t_to_slv(x : uint1908_t) return std_logic_vector;
function slv_to_uint1908_t(x : std_logic_vector) return uint1908_t;
subtype int1908_t is signed(1907 downto 0);
constant int1908_t_SLV_LEN : integer := 1908;
function int1908_t_to_slv(x : int1908_t) return std_logic_vector;
function slv_to_int1908_t(x : std_logic_vector) return int1908_t;
subtype uint1909_t is unsigned(1908 downto 0);
constant uint1909_t_SLV_LEN : integer := 1909;
function uint1909_t_to_slv(x : uint1909_t) return std_logic_vector;
function slv_to_uint1909_t(x : std_logic_vector) return uint1909_t;
subtype int1909_t is signed(1908 downto 0);
constant int1909_t_SLV_LEN : integer := 1909;
function int1909_t_to_slv(x : int1909_t) return std_logic_vector;
function slv_to_int1909_t(x : std_logic_vector) return int1909_t;
subtype uint1910_t is unsigned(1909 downto 0);
constant uint1910_t_SLV_LEN : integer := 1910;
function uint1910_t_to_slv(x : uint1910_t) return std_logic_vector;
function slv_to_uint1910_t(x : std_logic_vector) return uint1910_t;
subtype int1910_t is signed(1909 downto 0);
constant int1910_t_SLV_LEN : integer := 1910;
function int1910_t_to_slv(x : int1910_t) return std_logic_vector;
function slv_to_int1910_t(x : std_logic_vector) return int1910_t;
subtype uint1911_t is unsigned(1910 downto 0);
constant uint1911_t_SLV_LEN : integer := 1911;
function uint1911_t_to_slv(x : uint1911_t) return std_logic_vector;
function slv_to_uint1911_t(x : std_logic_vector) return uint1911_t;
subtype int1911_t is signed(1910 downto 0);
constant int1911_t_SLV_LEN : integer := 1911;
function int1911_t_to_slv(x : int1911_t) return std_logic_vector;
function slv_to_int1911_t(x : std_logic_vector) return int1911_t;
subtype uint1912_t is unsigned(1911 downto 0);
constant uint1912_t_SLV_LEN : integer := 1912;
function uint1912_t_to_slv(x : uint1912_t) return std_logic_vector;
function slv_to_uint1912_t(x : std_logic_vector) return uint1912_t;
subtype int1912_t is signed(1911 downto 0);
constant int1912_t_SLV_LEN : integer := 1912;
function int1912_t_to_slv(x : int1912_t) return std_logic_vector;
function slv_to_int1912_t(x : std_logic_vector) return int1912_t;
subtype uint1913_t is unsigned(1912 downto 0);
constant uint1913_t_SLV_LEN : integer := 1913;
function uint1913_t_to_slv(x : uint1913_t) return std_logic_vector;
function slv_to_uint1913_t(x : std_logic_vector) return uint1913_t;
subtype int1913_t is signed(1912 downto 0);
constant int1913_t_SLV_LEN : integer := 1913;
function int1913_t_to_slv(x : int1913_t) return std_logic_vector;
function slv_to_int1913_t(x : std_logic_vector) return int1913_t;
subtype uint1914_t is unsigned(1913 downto 0);
constant uint1914_t_SLV_LEN : integer := 1914;
function uint1914_t_to_slv(x : uint1914_t) return std_logic_vector;
function slv_to_uint1914_t(x : std_logic_vector) return uint1914_t;
subtype int1914_t is signed(1913 downto 0);
constant int1914_t_SLV_LEN : integer := 1914;
function int1914_t_to_slv(x : int1914_t) return std_logic_vector;
function slv_to_int1914_t(x : std_logic_vector) return int1914_t;
subtype uint1915_t is unsigned(1914 downto 0);
constant uint1915_t_SLV_LEN : integer := 1915;
function uint1915_t_to_slv(x : uint1915_t) return std_logic_vector;
function slv_to_uint1915_t(x : std_logic_vector) return uint1915_t;
subtype int1915_t is signed(1914 downto 0);
constant int1915_t_SLV_LEN : integer := 1915;
function int1915_t_to_slv(x : int1915_t) return std_logic_vector;
function slv_to_int1915_t(x : std_logic_vector) return int1915_t;
subtype uint1916_t is unsigned(1915 downto 0);
constant uint1916_t_SLV_LEN : integer := 1916;
function uint1916_t_to_slv(x : uint1916_t) return std_logic_vector;
function slv_to_uint1916_t(x : std_logic_vector) return uint1916_t;
subtype int1916_t is signed(1915 downto 0);
constant int1916_t_SLV_LEN : integer := 1916;
function int1916_t_to_slv(x : int1916_t) return std_logic_vector;
function slv_to_int1916_t(x : std_logic_vector) return int1916_t;
subtype uint1917_t is unsigned(1916 downto 0);
constant uint1917_t_SLV_LEN : integer := 1917;
function uint1917_t_to_slv(x : uint1917_t) return std_logic_vector;
function slv_to_uint1917_t(x : std_logic_vector) return uint1917_t;
subtype int1917_t is signed(1916 downto 0);
constant int1917_t_SLV_LEN : integer := 1917;
function int1917_t_to_slv(x : int1917_t) return std_logic_vector;
function slv_to_int1917_t(x : std_logic_vector) return int1917_t;
subtype uint1918_t is unsigned(1917 downto 0);
constant uint1918_t_SLV_LEN : integer := 1918;
function uint1918_t_to_slv(x : uint1918_t) return std_logic_vector;
function slv_to_uint1918_t(x : std_logic_vector) return uint1918_t;
subtype int1918_t is signed(1917 downto 0);
constant int1918_t_SLV_LEN : integer := 1918;
function int1918_t_to_slv(x : int1918_t) return std_logic_vector;
function slv_to_int1918_t(x : std_logic_vector) return int1918_t;
subtype uint1919_t is unsigned(1918 downto 0);
constant uint1919_t_SLV_LEN : integer := 1919;
function uint1919_t_to_slv(x : uint1919_t) return std_logic_vector;
function slv_to_uint1919_t(x : std_logic_vector) return uint1919_t;
subtype int1919_t is signed(1918 downto 0);
constant int1919_t_SLV_LEN : integer := 1919;
function int1919_t_to_slv(x : int1919_t) return std_logic_vector;
function slv_to_int1919_t(x : std_logic_vector) return int1919_t;
subtype uint1920_t is unsigned(1919 downto 0);
constant uint1920_t_SLV_LEN : integer := 1920;
function uint1920_t_to_slv(x : uint1920_t) return std_logic_vector;
function slv_to_uint1920_t(x : std_logic_vector) return uint1920_t;
subtype int1920_t is signed(1919 downto 0);
constant int1920_t_SLV_LEN : integer := 1920;
function int1920_t_to_slv(x : int1920_t) return std_logic_vector;
function slv_to_int1920_t(x : std_logic_vector) return int1920_t;
subtype uint1921_t is unsigned(1920 downto 0);
constant uint1921_t_SLV_LEN : integer := 1921;
function uint1921_t_to_slv(x : uint1921_t) return std_logic_vector;
function slv_to_uint1921_t(x : std_logic_vector) return uint1921_t;
subtype int1921_t is signed(1920 downto 0);
constant int1921_t_SLV_LEN : integer := 1921;
function int1921_t_to_slv(x : int1921_t) return std_logic_vector;
function slv_to_int1921_t(x : std_logic_vector) return int1921_t;
subtype uint1922_t is unsigned(1921 downto 0);
constant uint1922_t_SLV_LEN : integer := 1922;
function uint1922_t_to_slv(x : uint1922_t) return std_logic_vector;
function slv_to_uint1922_t(x : std_logic_vector) return uint1922_t;
subtype int1922_t is signed(1921 downto 0);
constant int1922_t_SLV_LEN : integer := 1922;
function int1922_t_to_slv(x : int1922_t) return std_logic_vector;
function slv_to_int1922_t(x : std_logic_vector) return int1922_t;
subtype uint1923_t is unsigned(1922 downto 0);
constant uint1923_t_SLV_LEN : integer := 1923;
function uint1923_t_to_slv(x : uint1923_t) return std_logic_vector;
function slv_to_uint1923_t(x : std_logic_vector) return uint1923_t;
subtype int1923_t is signed(1922 downto 0);
constant int1923_t_SLV_LEN : integer := 1923;
function int1923_t_to_slv(x : int1923_t) return std_logic_vector;
function slv_to_int1923_t(x : std_logic_vector) return int1923_t;
subtype uint1924_t is unsigned(1923 downto 0);
constant uint1924_t_SLV_LEN : integer := 1924;
function uint1924_t_to_slv(x : uint1924_t) return std_logic_vector;
function slv_to_uint1924_t(x : std_logic_vector) return uint1924_t;
subtype int1924_t is signed(1923 downto 0);
constant int1924_t_SLV_LEN : integer := 1924;
function int1924_t_to_slv(x : int1924_t) return std_logic_vector;
function slv_to_int1924_t(x : std_logic_vector) return int1924_t;
subtype uint1925_t is unsigned(1924 downto 0);
constant uint1925_t_SLV_LEN : integer := 1925;
function uint1925_t_to_slv(x : uint1925_t) return std_logic_vector;
function slv_to_uint1925_t(x : std_logic_vector) return uint1925_t;
subtype int1925_t is signed(1924 downto 0);
constant int1925_t_SLV_LEN : integer := 1925;
function int1925_t_to_slv(x : int1925_t) return std_logic_vector;
function slv_to_int1925_t(x : std_logic_vector) return int1925_t;
subtype uint1926_t is unsigned(1925 downto 0);
constant uint1926_t_SLV_LEN : integer := 1926;
function uint1926_t_to_slv(x : uint1926_t) return std_logic_vector;
function slv_to_uint1926_t(x : std_logic_vector) return uint1926_t;
subtype int1926_t is signed(1925 downto 0);
constant int1926_t_SLV_LEN : integer := 1926;
function int1926_t_to_slv(x : int1926_t) return std_logic_vector;
function slv_to_int1926_t(x : std_logic_vector) return int1926_t;
subtype uint1927_t is unsigned(1926 downto 0);
constant uint1927_t_SLV_LEN : integer := 1927;
function uint1927_t_to_slv(x : uint1927_t) return std_logic_vector;
function slv_to_uint1927_t(x : std_logic_vector) return uint1927_t;
subtype int1927_t is signed(1926 downto 0);
constant int1927_t_SLV_LEN : integer := 1927;
function int1927_t_to_slv(x : int1927_t) return std_logic_vector;
function slv_to_int1927_t(x : std_logic_vector) return int1927_t;
subtype uint1928_t is unsigned(1927 downto 0);
constant uint1928_t_SLV_LEN : integer := 1928;
function uint1928_t_to_slv(x : uint1928_t) return std_logic_vector;
function slv_to_uint1928_t(x : std_logic_vector) return uint1928_t;
subtype int1928_t is signed(1927 downto 0);
constant int1928_t_SLV_LEN : integer := 1928;
function int1928_t_to_slv(x : int1928_t) return std_logic_vector;
function slv_to_int1928_t(x : std_logic_vector) return int1928_t;
subtype uint1929_t is unsigned(1928 downto 0);
constant uint1929_t_SLV_LEN : integer := 1929;
function uint1929_t_to_slv(x : uint1929_t) return std_logic_vector;
function slv_to_uint1929_t(x : std_logic_vector) return uint1929_t;
subtype int1929_t is signed(1928 downto 0);
constant int1929_t_SLV_LEN : integer := 1929;
function int1929_t_to_slv(x : int1929_t) return std_logic_vector;
function slv_to_int1929_t(x : std_logic_vector) return int1929_t;
subtype uint1930_t is unsigned(1929 downto 0);
constant uint1930_t_SLV_LEN : integer := 1930;
function uint1930_t_to_slv(x : uint1930_t) return std_logic_vector;
function slv_to_uint1930_t(x : std_logic_vector) return uint1930_t;
subtype int1930_t is signed(1929 downto 0);
constant int1930_t_SLV_LEN : integer := 1930;
function int1930_t_to_slv(x : int1930_t) return std_logic_vector;
function slv_to_int1930_t(x : std_logic_vector) return int1930_t;
subtype uint1931_t is unsigned(1930 downto 0);
constant uint1931_t_SLV_LEN : integer := 1931;
function uint1931_t_to_slv(x : uint1931_t) return std_logic_vector;
function slv_to_uint1931_t(x : std_logic_vector) return uint1931_t;
subtype int1931_t is signed(1930 downto 0);
constant int1931_t_SLV_LEN : integer := 1931;
function int1931_t_to_slv(x : int1931_t) return std_logic_vector;
function slv_to_int1931_t(x : std_logic_vector) return int1931_t;
subtype uint1932_t is unsigned(1931 downto 0);
constant uint1932_t_SLV_LEN : integer := 1932;
function uint1932_t_to_slv(x : uint1932_t) return std_logic_vector;
function slv_to_uint1932_t(x : std_logic_vector) return uint1932_t;
subtype int1932_t is signed(1931 downto 0);
constant int1932_t_SLV_LEN : integer := 1932;
function int1932_t_to_slv(x : int1932_t) return std_logic_vector;
function slv_to_int1932_t(x : std_logic_vector) return int1932_t;
subtype uint1933_t is unsigned(1932 downto 0);
constant uint1933_t_SLV_LEN : integer := 1933;
function uint1933_t_to_slv(x : uint1933_t) return std_logic_vector;
function slv_to_uint1933_t(x : std_logic_vector) return uint1933_t;
subtype int1933_t is signed(1932 downto 0);
constant int1933_t_SLV_LEN : integer := 1933;
function int1933_t_to_slv(x : int1933_t) return std_logic_vector;
function slv_to_int1933_t(x : std_logic_vector) return int1933_t;
subtype uint1934_t is unsigned(1933 downto 0);
constant uint1934_t_SLV_LEN : integer := 1934;
function uint1934_t_to_slv(x : uint1934_t) return std_logic_vector;
function slv_to_uint1934_t(x : std_logic_vector) return uint1934_t;
subtype int1934_t is signed(1933 downto 0);
constant int1934_t_SLV_LEN : integer := 1934;
function int1934_t_to_slv(x : int1934_t) return std_logic_vector;
function slv_to_int1934_t(x : std_logic_vector) return int1934_t;
subtype uint1935_t is unsigned(1934 downto 0);
constant uint1935_t_SLV_LEN : integer := 1935;
function uint1935_t_to_slv(x : uint1935_t) return std_logic_vector;
function slv_to_uint1935_t(x : std_logic_vector) return uint1935_t;
subtype int1935_t is signed(1934 downto 0);
constant int1935_t_SLV_LEN : integer := 1935;
function int1935_t_to_slv(x : int1935_t) return std_logic_vector;
function slv_to_int1935_t(x : std_logic_vector) return int1935_t;
subtype uint1936_t is unsigned(1935 downto 0);
constant uint1936_t_SLV_LEN : integer := 1936;
function uint1936_t_to_slv(x : uint1936_t) return std_logic_vector;
function slv_to_uint1936_t(x : std_logic_vector) return uint1936_t;
subtype int1936_t is signed(1935 downto 0);
constant int1936_t_SLV_LEN : integer := 1936;
function int1936_t_to_slv(x : int1936_t) return std_logic_vector;
function slv_to_int1936_t(x : std_logic_vector) return int1936_t;
subtype uint1937_t is unsigned(1936 downto 0);
constant uint1937_t_SLV_LEN : integer := 1937;
function uint1937_t_to_slv(x : uint1937_t) return std_logic_vector;
function slv_to_uint1937_t(x : std_logic_vector) return uint1937_t;
subtype int1937_t is signed(1936 downto 0);
constant int1937_t_SLV_LEN : integer := 1937;
function int1937_t_to_slv(x : int1937_t) return std_logic_vector;
function slv_to_int1937_t(x : std_logic_vector) return int1937_t;
subtype uint1938_t is unsigned(1937 downto 0);
constant uint1938_t_SLV_LEN : integer := 1938;
function uint1938_t_to_slv(x : uint1938_t) return std_logic_vector;
function slv_to_uint1938_t(x : std_logic_vector) return uint1938_t;
subtype int1938_t is signed(1937 downto 0);
constant int1938_t_SLV_LEN : integer := 1938;
function int1938_t_to_slv(x : int1938_t) return std_logic_vector;
function slv_to_int1938_t(x : std_logic_vector) return int1938_t;
subtype uint1939_t is unsigned(1938 downto 0);
constant uint1939_t_SLV_LEN : integer := 1939;
function uint1939_t_to_slv(x : uint1939_t) return std_logic_vector;
function slv_to_uint1939_t(x : std_logic_vector) return uint1939_t;
subtype int1939_t is signed(1938 downto 0);
constant int1939_t_SLV_LEN : integer := 1939;
function int1939_t_to_slv(x : int1939_t) return std_logic_vector;
function slv_to_int1939_t(x : std_logic_vector) return int1939_t;
subtype uint1940_t is unsigned(1939 downto 0);
constant uint1940_t_SLV_LEN : integer := 1940;
function uint1940_t_to_slv(x : uint1940_t) return std_logic_vector;
function slv_to_uint1940_t(x : std_logic_vector) return uint1940_t;
subtype int1940_t is signed(1939 downto 0);
constant int1940_t_SLV_LEN : integer := 1940;
function int1940_t_to_slv(x : int1940_t) return std_logic_vector;
function slv_to_int1940_t(x : std_logic_vector) return int1940_t;
subtype uint1941_t is unsigned(1940 downto 0);
constant uint1941_t_SLV_LEN : integer := 1941;
function uint1941_t_to_slv(x : uint1941_t) return std_logic_vector;
function slv_to_uint1941_t(x : std_logic_vector) return uint1941_t;
subtype int1941_t is signed(1940 downto 0);
constant int1941_t_SLV_LEN : integer := 1941;
function int1941_t_to_slv(x : int1941_t) return std_logic_vector;
function slv_to_int1941_t(x : std_logic_vector) return int1941_t;
subtype uint1942_t is unsigned(1941 downto 0);
constant uint1942_t_SLV_LEN : integer := 1942;
function uint1942_t_to_slv(x : uint1942_t) return std_logic_vector;
function slv_to_uint1942_t(x : std_logic_vector) return uint1942_t;
subtype int1942_t is signed(1941 downto 0);
constant int1942_t_SLV_LEN : integer := 1942;
function int1942_t_to_slv(x : int1942_t) return std_logic_vector;
function slv_to_int1942_t(x : std_logic_vector) return int1942_t;
subtype uint1943_t is unsigned(1942 downto 0);
constant uint1943_t_SLV_LEN : integer := 1943;
function uint1943_t_to_slv(x : uint1943_t) return std_logic_vector;
function slv_to_uint1943_t(x : std_logic_vector) return uint1943_t;
subtype int1943_t is signed(1942 downto 0);
constant int1943_t_SLV_LEN : integer := 1943;
function int1943_t_to_slv(x : int1943_t) return std_logic_vector;
function slv_to_int1943_t(x : std_logic_vector) return int1943_t;
subtype uint1944_t is unsigned(1943 downto 0);
constant uint1944_t_SLV_LEN : integer := 1944;
function uint1944_t_to_slv(x : uint1944_t) return std_logic_vector;
function slv_to_uint1944_t(x : std_logic_vector) return uint1944_t;
subtype int1944_t is signed(1943 downto 0);
constant int1944_t_SLV_LEN : integer := 1944;
function int1944_t_to_slv(x : int1944_t) return std_logic_vector;
function slv_to_int1944_t(x : std_logic_vector) return int1944_t;
subtype uint1945_t is unsigned(1944 downto 0);
constant uint1945_t_SLV_LEN : integer := 1945;
function uint1945_t_to_slv(x : uint1945_t) return std_logic_vector;
function slv_to_uint1945_t(x : std_logic_vector) return uint1945_t;
subtype int1945_t is signed(1944 downto 0);
constant int1945_t_SLV_LEN : integer := 1945;
function int1945_t_to_slv(x : int1945_t) return std_logic_vector;
function slv_to_int1945_t(x : std_logic_vector) return int1945_t;
subtype uint1946_t is unsigned(1945 downto 0);
constant uint1946_t_SLV_LEN : integer := 1946;
function uint1946_t_to_slv(x : uint1946_t) return std_logic_vector;
function slv_to_uint1946_t(x : std_logic_vector) return uint1946_t;
subtype int1946_t is signed(1945 downto 0);
constant int1946_t_SLV_LEN : integer := 1946;
function int1946_t_to_slv(x : int1946_t) return std_logic_vector;
function slv_to_int1946_t(x : std_logic_vector) return int1946_t;
subtype uint1947_t is unsigned(1946 downto 0);
constant uint1947_t_SLV_LEN : integer := 1947;
function uint1947_t_to_slv(x : uint1947_t) return std_logic_vector;
function slv_to_uint1947_t(x : std_logic_vector) return uint1947_t;
subtype int1947_t is signed(1946 downto 0);
constant int1947_t_SLV_LEN : integer := 1947;
function int1947_t_to_slv(x : int1947_t) return std_logic_vector;
function slv_to_int1947_t(x : std_logic_vector) return int1947_t;
subtype uint1948_t is unsigned(1947 downto 0);
constant uint1948_t_SLV_LEN : integer := 1948;
function uint1948_t_to_slv(x : uint1948_t) return std_logic_vector;
function slv_to_uint1948_t(x : std_logic_vector) return uint1948_t;
subtype int1948_t is signed(1947 downto 0);
constant int1948_t_SLV_LEN : integer := 1948;
function int1948_t_to_slv(x : int1948_t) return std_logic_vector;
function slv_to_int1948_t(x : std_logic_vector) return int1948_t;
subtype uint1949_t is unsigned(1948 downto 0);
constant uint1949_t_SLV_LEN : integer := 1949;
function uint1949_t_to_slv(x : uint1949_t) return std_logic_vector;
function slv_to_uint1949_t(x : std_logic_vector) return uint1949_t;
subtype int1949_t is signed(1948 downto 0);
constant int1949_t_SLV_LEN : integer := 1949;
function int1949_t_to_slv(x : int1949_t) return std_logic_vector;
function slv_to_int1949_t(x : std_logic_vector) return int1949_t;
subtype uint1950_t is unsigned(1949 downto 0);
constant uint1950_t_SLV_LEN : integer := 1950;
function uint1950_t_to_slv(x : uint1950_t) return std_logic_vector;
function slv_to_uint1950_t(x : std_logic_vector) return uint1950_t;
subtype int1950_t is signed(1949 downto 0);
constant int1950_t_SLV_LEN : integer := 1950;
function int1950_t_to_slv(x : int1950_t) return std_logic_vector;
function slv_to_int1950_t(x : std_logic_vector) return int1950_t;
subtype uint1951_t is unsigned(1950 downto 0);
constant uint1951_t_SLV_LEN : integer := 1951;
function uint1951_t_to_slv(x : uint1951_t) return std_logic_vector;
function slv_to_uint1951_t(x : std_logic_vector) return uint1951_t;
subtype int1951_t is signed(1950 downto 0);
constant int1951_t_SLV_LEN : integer := 1951;
function int1951_t_to_slv(x : int1951_t) return std_logic_vector;
function slv_to_int1951_t(x : std_logic_vector) return int1951_t;
subtype uint1952_t is unsigned(1951 downto 0);
constant uint1952_t_SLV_LEN : integer := 1952;
function uint1952_t_to_slv(x : uint1952_t) return std_logic_vector;
function slv_to_uint1952_t(x : std_logic_vector) return uint1952_t;
subtype int1952_t is signed(1951 downto 0);
constant int1952_t_SLV_LEN : integer := 1952;
function int1952_t_to_slv(x : int1952_t) return std_logic_vector;
function slv_to_int1952_t(x : std_logic_vector) return int1952_t;
subtype uint1953_t is unsigned(1952 downto 0);
constant uint1953_t_SLV_LEN : integer := 1953;
function uint1953_t_to_slv(x : uint1953_t) return std_logic_vector;
function slv_to_uint1953_t(x : std_logic_vector) return uint1953_t;
subtype int1953_t is signed(1952 downto 0);
constant int1953_t_SLV_LEN : integer := 1953;
function int1953_t_to_slv(x : int1953_t) return std_logic_vector;
function slv_to_int1953_t(x : std_logic_vector) return int1953_t;
subtype uint1954_t is unsigned(1953 downto 0);
constant uint1954_t_SLV_LEN : integer := 1954;
function uint1954_t_to_slv(x : uint1954_t) return std_logic_vector;
function slv_to_uint1954_t(x : std_logic_vector) return uint1954_t;
subtype int1954_t is signed(1953 downto 0);
constant int1954_t_SLV_LEN : integer := 1954;
function int1954_t_to_slv(x : int1954_t) return std_logic_vector;
function slv_to_int1954_t(x : std_logic_vector) return int1954_t;
subtype uint1955_t is unsigned(1954 downto 0);
constant uint1955_t_SLV_LEN : integer := 1955;
function uint1955_t_to_slv(x : uint1955_t) return std_logic_vector;
function slv_to_uint1955_t(x : std_logic_vector) return uint1955_t;
subtype int1955_t is signed(1954 downto 0);
constant int1955_t_SLV_LEN : integer := 1955;
function int1955_t_to_slv(x : int1955_t) return std_logic_vector;
function slv_to_int1955_t(x : std_logic_vector) return int1955_t;
subtype uint1956_t is unsigned(1955 downto 0);
constant uint1956_t_SLV_LEN : integer := 1956;
function uint1956_t_to_slv(x : uint1956_t) return std_logic_vector;
function slv_to_uint1956_t(x : std_logic_vector) return uint1956_t;
subtype int1956_t is signed(1955 downto 0);
constant int1956_t_SLV_LEN : integer := 1956;
function int1956_t_to_slv(x : int1956_t) return std_logic_vector;
function slv_to_int1956_t(x : std_logic_vector) return int1956_t;
subtype uint1957_t is unsigned(1956 downto 0);
constant uint1957_t_SLV_LEN : integer := 1957;
function uint1957_t_to_slv(x : uint1957_t) return std_logic_vector;
function slv_to_uint1957_t(x : std_logic_vector) return uint1957_t;
subtype int1957_t is signed(1956 downto 0);
constant int1957_t_SLV_LEN : integer := 1957;
function int1957_t_to_slv(x : int1957_t) return std_logic_vector;
function slv_to_int1957_t(x : std_logic_vector) return int1957_t;
subtype uint1958_t is unsigned(1957 downto 0);
constant uint1958_t_SLV_LEN : integer := 1958;
function uint1958_t_to_slv(x : uint1958_t) return std_logic_vector;
function slv_to_uint1958_t(x : std_logic_vector) return uint1958_t;
subtype int1958_t is signed(1957 downto 0);
constant int1958_t_SLV_LEN : integer := 1958;
function int1958_t_to_slv(x : int1958_t) return std_logic_vector;
function slv_to_int1958_t(x : std_logic_vector) return int1958_t;
subtype uint1959_t is unsigned(1958 downto 0);
constant uint1959_t_SLV_LEN : integer := 1959;
function uint1959_t_to_slv(x : uint1959_t) return std_logic_vector;
function slv_to_uint1959_t(x : std_logic_vector) return uint1959_t;
subtype int1959_t is signed(1958 downto 0);
constant int1959_t_SLV_LEN : integer := 1959;
function int1959_t_to_slv(x : int1959_t) return std_logic_vector;
function slv_to_int1959_t(x : std_logic_vector) return int1959_t;
subtype uint1960_t is unsigned(1959 downto 0);
constant uint1960_t_SLV_LEN : integer := 1960;
function uint1960_t_to_slv(x : uint1960_t) return std_logic_vector;
function slv_to_uint1960_t(x : std_logic_vector) return uint1960_t;
subtype int1960_t is signed(1959 downto 0);
constant int1960_t_SLV_LEN : integer := 1960;
function int1960_t_to_slv(x : int1960_t) return std_logic_vector;
function slv_to_int1960_t(x : std_logic_vector) return int1960_t;
subtype uint1961_t is unsigned(1960 downto 0);
constant uint1961_t_SLV_LEN : integer := 1961;
function uint1961_t_to_slv(x : uint1961_t) return std_logic_vector;
function slv_to_uint1961_t(x : std_logic_vector) return uint1961_t;
subtype int1961_t is signed(1960 downto 0);
constant int1961_t_SLV_LEN : integer := 1961;
function int1961_t_to_slv(x : int1961_t) return std_logic_vector;
function slv_to_int1961_t(x : std_logic_vector) return int1961_t;
subtype uint1962_t is unsigned(1961 downto 0);
constant uint1962_t_SLV_LEN : integer := 1962;
function uint1962_t_to_slv(x : uint1962_t) return std_logic_vector;
function slv_to_uint1962_t(x : std_logic_vector) return uint1962_t;
subtype int1962_t is signed(1961 downto 0);
constant int1962_t_SLV_LEN : integer := 1962;
function int1962_t_to_slv(x : int1962_t) return std_logic_vector;
function slv_to_int1962_t(x : std_logic_vector) return int1962_t;
subtype uint1963_t is unsigned(1962 downto 0);
constant uint1963_t_SLV_LEN : integer := 1963;
function uint1963_t_to_slv(x : uint1963_t) return std_logic_vector;
function slv_to_uint1963_t(x : std_logic_vector) return uint1963_t;
subtype int1963_t is signed(1962 downto 0);
constant int1963_t_SLV_LEN : integer := 1963;
function int1963_t_to_slv(x : int1963_t) return std_logic_vector;
function slv_to_int1963_t(x : std_logic_vector) return int1963_t;
subtype uint1964_t is unsigned(1963 downto 0);
constant uint1964_t_SLV_LEN : integer := 1964;
function uint1964_t_to_slv(x : uint1964_t) return std_logic_vector;
function slv_to_uint1964_t(x : std_logic_vector) return uint1964_t;
subtype int1964_t is signed(1963 downto 0);
constant int1964_t_SLV_LEN : integer := 1964;
function int1964_t_to_slv(x : int1964_t) return std_logic_vector;
function slv_to_int1964_t(x : std_logic_vector) return int1964_t;
subtype uint1965_t is unsigned(1964 downto 0);
constant uint1965_t_SLV_LEN : integer := 1965;
function uint1965_t_to_slv(x : uint1965_t) return std_logic_vector;
function slv_to_uint1965_t(x : std_logic_vector) return uint1965_t;
subtype int1965_t is signed(1964 downto 0);
constant int1965_t_SLV_LEN : integer := 1965;
function int1965_t_to_slv(x : int1965_t) return std_logic_vector;
function slv_to_int1965_t(x : std_logic_vector) return int1965_t;
subtype uint1966_t is unsigned(1965 downto 0);
constant uint1966_t_SLV_LEN : integer := 1966;
function uint1966_t_to_slv(x : uint1966_t) return std_logic_vector;
function slv_to_uint1966_t(x : std_logic_vector) return uint1966_t;
subtype int1966_t is signed(1965 downto 0);
constant int1966_t_SLV_LEN : integer := 1966;
function int1966_t_to_slv(x : int1966_t) return std_logic_vector;
function slv_to_int1966_t(x : std_logic_vector) return int1966_t;
subtype uint1967_t is unsigned(1966 downto 0);
constant uint1967_t_SLV_LEN : integer := 1967;
function uint1967_t_to_slv(x : uint1967_t) return std_logic_vector;
function slv_to_uint1967_t(x : std_logic_vector) return uint1967_t;
subtype int1967_t is signed(1966 downto 0);
constant int1967_t_SLV_LEN : integer := 1967;
function int1967_t_to_slv(x : int1967_t) return std_logic_vector;
function slv_to_int1967_t(x : std_logic_vector) return int1967_t;
subtype uint1968_t is unsigned(1967 downto 0);
constant uint1968_t_SLV_LEN : integer := 1968;
function uint1968_t_to_slv(x : uint1968_t) return std_logic_vector;
function slv_to_uint1968_t(x : std_logic_vector) return uint1968_t;
subtype int1968_t is signed(1967 downto 0);
constant int1968_t_SLV_LEN : integer := 1968;
function int1968_t_to_slv(x : int1968_t) return std_logic_vector;
function slv_to_int1968_t(x : std_logic_vector) return int1968_t;
subtype uint1969_t is unsigned(1968 downto 0);
constant uint1969_t_SLV_LEN : integer := 1969;
function uint1969_t_to_slv(x : uint1969_t) return std_logic_vector;
function slv_to_uint1969_t(x : std_logic_vector) return uint1969_t;
subtype int1969_t is signed(1968 downto 0);
constant int1969_t_SLV_LEN : integer := 1969;
function int1969_t_to_slv(x : int1969_t) return std_logic_vector;
function slv_to_int1969_t(x : std_logic_vector) return int1969_t;
subtype uint1970_t is unsigned(1969 downto 0);
constant uint1970_t_SLV_LEN : integer := 1970;
function uint1970_t_to_slv(x : uint1970_t) return std_logic_vector;
function slv_to_uint1970_t(x : std_logic_vector) return uint1970_t;
subtype int1970_t is signed(1969 downto 0);
constant int1970_t_SLV_LEN : integer := 1970;
function int1970_t_to_slv(x : int1970_t) return std_logic_vector;
function slv_to_int1970_t(x : std_logic_vector) return int1970_t;
subtype uint1971_t is unsigned(1970 downto 0);
constant uint1971_t_SLV_LEN : integer := 1971;
function uint1971_t_to_slv(x : uint1971_t) return std_logic_vector;
function slv_to_uint1971_t(x : std_logic_vector) return uint1971_t;
subtype int1971_t is signed(1970 downto 0);
constant int1971_t_SLV_LEN : integer := 1971;
function int1971_t_to_slv(x : int1971_t) return std_logic_vector;
function slv_to_int1971_t(x : std_logic_vector) return int1971_t;
subtype uint1972_t is unsigned(1971 downto 0);
constant uint1972_t_SLV_LEN : integer := 1972;
function uint1972_t_to_slv(x : uint1972_t) return std_logic_vector;
function slv_to_uint1972_t(x : std_logic_vector) return uint1972_t;
subtype int1972_t is signed(1971 downto 0);
constant int1972_t_SLV_LEN : integer := 1972;
function int1972_t_to_slv(x : int1972_t) return std_logic_vector;
function slv_to_int1972_t(x : std_logic_vector) return int1972_t;
subtype uint1973_t is unsigned(1972 downto 0);
constant uint1973_t_SLV_LEN : integer := 1973;
function uint1973_t_to_slv(x : uint1973_t) return std_logic_vector;
function slv_to_uint1973_t(x : std_logic_vector) return uint1973_t;
subtype int1973_t is signed(1972 downto 0);
constant int1973_t_SLV_LEN : integer := 1973;
function int1973_t_to_slv(x : int1973_t) return std_logic_vector;
function slv_to_int1973_t(x : std_logic_vector) return int1973_t;
subtype uint1974_t is unsigned(1973 downto 0);
constant uint1974_t_SLV_LEN : integer := 1974;
function uint1974_t_to_slv(x : uint1974_t) return std_logic_vector;
function slv_to_uint1974_t(x : std_logic_vector) return uint1974_t;
subtype int1974_t is signed(1973 downto 0);
constant int1974_t_SLV_LEN : integer := 1974;
function int1974_t_to_slv(x : int1974_t) return std_logic_vector;
function slv_to_int1974_t(x : std_logic_vector) return int1974_t;
subtype uint1975_t is unsigned(1974 downto 0);
constant uint1975_t_SLV_LEN : integer := 1975;
function uint1975_t_to_slv(x : uint1975_t) return std_logic_vector;
function slv_to_uint1975_t(x : std_logic_vector) return uint1975_t;
subtype int1975_t is signed(1974 downto 0);
constant int1975_t_SLV_LEN : integer := 1975;
function int1975_t_to_slv(x : int1975_t) return std_logic_vector;
function slv_to_int1975_t(x : std_logic_vector) return int1975_t;
subtype uint1976_t is unsigned(1975 downto 0);
constant uint1976_t_SLV_LEN : integer := 1976;
function uint1976_t_to_slv(x : uint1976_t) return std_logic_vector;
function slv_to_uint1976_t(x : std_logic_vector) return uint1976_t;
subtype int1976_t is signed(1975 downto 0);
constant int1976_t_SLV_LEN : integer := 1976;
function int1976_t_to_slv(x : int1976_t) return std_logic_vector;
function slv_to_int1976_t(x : std_logic_vector) return int1976_t;
subtype uint1977_t is unsigned(1976 downto 0);
constant uint1977_t_SLV_LEN : integer := 1977;
function uint1977_t_to_slv(x : uint1977_t) return std_logic_vector;
function slv_to_uint1977_t(x : std_logic_vector) return uint1977_t;
subtype int1977_t is signed(1976 downto 0);
constant int1977_t_SLV_LEN : integer := 1977;
function int1977_t_to_slv(x : int1977_t) return std_logic_vector;
function slv_to_int1977_t(x : std_logic_vector) return int1977_t;
subtype uint1978_t is unsigned(1977 downto 0);
constant uint1978_t_SLV_LEN : integer := 1978;
function uint1978_t_to_slv(x : uint1978_t) return std_logic_vector;
function slv_to_uint1978_t(x : std_logic_vector) return uint1978_t;
subtype int1978_t is signed(1977 downto 0);
constant int1978_t_SLV_LEN : integer := 1978;
function int1978_t_to_slv(x : int1978_t) return std_logic_vector;
function slv_to_int1978_t(x : std_logic_vector) return int1978_t;
subtype uint1979_t is unsigned(1978 downto 0);
constant uint1979_t_SLV_LEN : integer := 1979;
function uint1979_t_to_slv(x : uint1979_t) return std_logic_vector;
function slv_to_uint1979_t(x : std_logic_vector) return uint1979_t;
subtype int1979_t is signed(1978 downto 0);
constant int1979_t_SLV_LEN : integer := 1979;
function int1979_t_to_slv(x : int1979_t) return std_logic_vector;
function slv_to_int1979_t(x : std_logic_vector) return int1979_t;
subtype uint1980_t is unsigned(1979 downto 0);
constant uint1980_t_SLV_LEN : integer := 1980;
function uint1980_t_to_slv(x : uint1980_t) return std_logic_vector;
function slv_to_uint1980_t(x : std_logic_vector) return uint1980_t;
subtype int1980_t is signed(1979 downto 0);
constant int1980_t_SLV_LEN : integer := 1980;
function int1980_t_to_slv(x : int1980_t) return std_logic_vector;
function slv_to_int1980_t(x : std_logic_vector) return int1980_t;
subtype uint1981_t is unsigned(1980 downto 0);
constant uint1981_t_SLV_LEN : integer := 1981;
function uint1981_t_to_slv(x : uint1981_t) return std_logic_vector;
function slv_to_uint1981_t(x : std_logic_vector) return uint1981_t;
subtype int1981_t is signed(1980 downto 0);
constant int1981_t_SLV_LEN : integer := 1981;
function int1981_t_to_slv(x : int1981_t) return std_logic_vector;
function slv_to_int1981_t(x : std_logic_vector) return int1981_t;
subtype uint1982_t is unsigned(1981 downto 0);
constant uint1982_t_SLV_LEN : integer := 1982;
function uint1982_t_to_slv(x : uint1982_t) return std_logic_vector;
function slv_to_uint1982_t(x : std_logic_vector) return uint1982_t;
subtype int1982_t is signed(1981 downto 0);
constant int1982_t_SLV_LEN : integer := 1982;
function int1982_t_to_slv(x : int1982_t) return std_logic_vector;
function slv_to_int1982_t(x : std_logic_vector) return int1982_t;
subtype uint1983_t is unsigned(1982 downto 0);
constant uint1983_t_SLV_LEN : integer := 1983;
function uint1983_t_to_slv(x : uint1983_t) return std_logic_vector;
function slv_to_uint1983_t(x : std_logic_vector) return uint1983_t;
subtype int1983_t is signed(1982 downto 0);
constant int1983_t_SLV_LEN : integer := 1983;
function int1983_t_to_slv(x : int1983_t) return std_logic_vector;
function slv_to_int1983_t(x : std_logic_vector) return int1983_t;
subtype uint1984_t is unsigned(1983 downto 0);
constant uint1984_t_SLV_LEN : integer := 1984;
function uint1984_t_to_slv(x : uint1984_t) return std_logic_vector;
function slv_to_uint1984_t(x : std_logic_vector) return uint1984_t;
subtype int1984_t is signed(1983 downto 0);
constant int1984_t_SLV_LEN : integer := 1984;
function int1984_t_to_slv(x : int1984_t) return std_logic_vector;
function slv_to_int1984_t(x : std_logic_vector) return int1984_t;
subtype uint1985_t is unsigned(1984 downto 0);
constant uint1985_t_SLV_LEN : integer := 1985;
function uint1985_t_to_slv(x : uint1985_t) return std_logic_vector;
function slv_to_uint1985_t(x : std_logic_vector) return uint1985_t;
subtype int1985_t is signed(1984 downto 0);
constant int1985_t_SLV_LEN : integer := 1985;
function int1985_t_to_slv(x : int1985_t) return std_logic_vector;
function slv_to_int1985_t(x : std_logic_vector) return int1985_t;
subtype uint1986_t is unsigned(1985 downto 0);
constant uint1986_t_SLV_LEN : integer := 1986;
function uint1986_t_to_slv(x : uint1986_t) return std_logic_vector;
function slv_to_uint1986_t(x : std_logic_vector) return uint1986_t;
subtype int1986_t is signed(1985 downto 0);
constant int1986_t_SLV_LEN : integer := 1986;
function int1986_t_to_slv(x : int1986_t) return std_logic_vector;
function slv_to_int1986_t(x : std_logic_vector) return int1986_t;
subtype uint1987_t is unsigned(1986 downto 0);
constant uint1987_t_SLV_LEN : integer := 1987;
function uint1987_t_to_slv(x : uint1987_t) return std_logic_vector;
function slv_to_uint1987_t(x : std_logic_vector) return uint1987_t;
subtype int1987_t is signed(1986 downto 0);
constant int1987_t_SLV_LEN : integer := 1987;
function int1987_t_to_slv(x : int1987_t) return std_logic_vector;
function slv_to_int1987_t(x : std_logic_vector) return int1987_t;
subtype uint1988_t is unsigned(1987 downto 0);
constant uint1988_t_SLV_LEN : integer := 1988;
function uint1988_t_to_slv(x : uint1988_t) return std_logic_vector;
function slv_to_uint1988_t(x : std_logic_vector) return uint1988_t;
subtype int1988_t is signed(1987 downto 0);
constant int1988_t_SLV_LEN : integer := 1988;
function int1988_t_to_slv(x : int1988_t) return std_logic_vector;
function slv_to_int1988_t(x : std_logic_vector) return int1988_t;
subtype uint1989_t is unsigned(1988 downto 0);
constant uint1989_t_SLV_LEN : integer := 1989;
function uint1989_t_to_slv(x : uint1989_t) return std_logic_vector;
function slv_to_uint1989_t(x : std_logic_vector) return uint1989_t;
subtype int1989_t is signed(1988 downto 0);
constant int1989_t_SLV_LEN : integer := 1989;
function int1989_t_to_slv(x : int1989_t) return std_logic_vector;
function slv_to_int1989_t(x : std_logic_vector) return int1989_t;
subtype uint1990_t is unsigned(1989 downto 0);
constant uint1990_t_SLV_LEN : integer := 1990;
function uint1990_t_to_slv(x : uint1990_t) return std_logic_vector;
function slv_to_uint1990_t(x : std_logic_vector) return uint1990_t;
subtype int1990_t is signed(1989 downto 0);
constant int1990_t_SLV_LEN : integer := 1990;
function int1990_t_to_slv(x : int1990_t) return std_logic_vector;
function slv_to_int1990_t(x : std_logic_vector) return int1990_t;
subtype uint1991_t is unsigned(1990 downto 0);
constant uint1991_t_SLV_LEN : integer := 1991;
function uint1991_t_to_slv(x : uint1991_t) return std_logic_vector;
function slv_to_uint1991_t(x : std_logic_vector) return uint1991_t;
subtype int1991_t is signed(1990 downto 0);
constant int1991_t_SLV_LEN : integer := 1991;
function int1991_t_to_slv(x : int1991_t) return std_logic_vector;
function slv_to_int1991_t(x : std_logic_vector) return int1991_t;
subtype uint1992_t is unsigned(1991 downto 0);
constant uint1992_t_SLV_LEN : integer := 1992;
function uint1992_t_to_slv(x : uint1992_t) return std_logic_vector;
function slv_to_uint1992_t(x : std_logic_vector) return uint1992_t;
subtype int1992_t is signed(1991 downto 0);
constant int1992_t_SLV_LEN : integer := 1992;
function int1992_t_to_slv(x : int1992_t) return std_logic_vector;
function slv_to_int1992_t(x : std_logic_vector) return int1992_t;
subtype uint1993_t is unsigned(1992 downto 0);
constant uint1993_t_SLV_LEN : integer := 1993;
function uint1993_t_to_slv(x : uint1993_t) return std_logic_vector;
function slv_to_uint1993_t(x : std_logic_vector) return uint1993_t;
subtype int1993_t is signed(1992 downto 0);
constant int1993_t_SLV_LEN : integer := 1993;
function int1993_t_to_slv(x : int1993_t) return std_logic_vector;
function slv_to_int1993_t(x : std_logic_vector) return int1993_t;
subtype uint1994_t is unsigned(1993 downto 0);
constant uint1994_t_SLV_LEN : integer := 1994;
function uint1994_t_to_slv(x : uint1994_t) return std_logic_vector;
function slv_to_uint1994_t(x : std_logic_vector) return uint1994_t;
subtype int1994_t is signed(1993 downto 0);
constant int1994_t_SLV_LEN : integer := 1994;
function int1994_t_to_slv(x : int1994_t) return std_logic_vector;
function slv_to_int1994_t(x : std_logic_vector) return int1994_t;
subtype uint1995_t is unsigned(1994 downto 0);
constant uint1995_t_SLV_LEN : integer := 1995;
function uint1995_t_to_slv(x : uint1995_t) return std_logic_vector;
function slv_to_uint1995_t(x : std_logic_vector) return uint1995_t;
subtype int1995_t is signed(1994 downto 0);
constant int1995_t_SLV_LEN : integer := 1995;
function int1995_t_to_slv(x : int1995_t) return std_logic_vector;
function slv_to_int1995_t(x : std_logic_vector) return int1995_t;
subtype uint1996_t is unsigned(1995 downto 0);
constant uint1996_t_SLV_LEN : integer := 1996;
function uint1996_t_to_slv(x : uint1996_t) return std_logic_vector;
function slv_to_uint1996_t(x : std_logic_vector) return uint1996_t;
subtype int1996_t is signed(1995 downto 0);
constant int1996_t_SLV_LEN : integer := 1996;
function int1996_t_to_slv(x : int1996_t) return std_logic_vector;
function slv_to_int1996_t(x : std_logic_vector) return int1996_t;
subtype uint1997_t is unsigned(1996 downto 0);
constant uint1997_t_SLV_LEN : integer := 1997;
function uint1997_t_to_slv(x : uint1997_t) return std_logic_vector;
function slv_to_uint1997_t(x : std_logic_vector) return uint1997_t;
subtype int1997_t is signed(1996 downto 0);
constant int1997_t_SLV_LEN : integer := 1997;
function int1997_t_to_slv(x : int1997_t) return std_logic_vector;
function slv_to_int1997_t(x : std_logic_vector) return int1997_t;
subtype uint1998_t is unsigned(1997 downto 0);
constant uint1998_t_SLV_LEN : integer := 1998;
function uint1998_t_to_slv(x : uint1998_t) return std_logic_vector;
function slv_to_uint1998_t(x : std_logic_vector) return uint1998_t;
subtype int1998_t is signed(1997 downto 0);
constant int1998_t_SLV_LEN : integer := 1998;
function int1998_t_to_slv(x : int1998_t) return std_logic_vector;
function slv_to_int1998_t(x : std_logic_vector) return int1998_t;
subtype uint1999_t is unsigned(1998 downto 0);
constant uint1999_t_SLV_LEN : integer := 1999;
function uint1999_t_to_slv(x : uint1999_t) return std_logic_vector;
function slv_to_uint1999_t(x : std_logic_vector) return uint1999_t;
subtype int1999_t is signed(1998 downto 0);
constant int1999_t_SLV_LEN : integer := 1999;
function int1999_t_to_slv(x : int1999_t) return std_logic_vector;
function slv_to_int1999_t(x : std_logic_vector) return int1999_t;
subtype uint2000_t is unsigned(1999 downto 0);
constant uint2000_t_SLV_LEN : integer := 2000;
function uint2000_t_to_slv(x : uint2000_t) return std_logic_vector;
function slv_to_uint2000_t(x : std_logic_vector) return uint2000_t;
subtype int2000_t is signed(1999 downto 0);
constant int2000_t_SLV_LEN : integer := 2000;
function int2000_t_to_slv(x : int2000_t) return std_logic_vector;
function slv_to_int2000_t(x : std_logic_vector) return int2000_t;
subtype uint2001_t is unsigned(2000 downto 0);
constant uint2001_t_SLV_LEN : integer := 2001;
function uint2001_t_to_slv(x : uint2001_t) return std_logic_vector;
function slv_to_uint2001_t(x : std_logic_vector) return uint2001_t;
subtype int2001_t is signed(2000 downto 0);
constant int2001_t_SLV_LEN : integer := 2001;
function int2001_t_to_slv(x : int2001_t) return std_logic_vector;
function slv_to_int2001_t(x : std_logic_vector) return int2001_t;
subtype uint2002_t is unsigned(2001 downto 0);
constant uint2002_t_SLV_LEN : integer := 2002;
function uint2002_t_to_slv(x : uint2002_t) return std_logic_vector;
function slv_to_uint2002_t(x : std_logic_vector) return uint2002_t;
subtype int2002_t is signed(2001 downto 0);
constant int2002_t_SLV_LEN : integer := 2002;
function int2002_t_to_slv(x : int2002_t) return std_logic_vector;
function slv_to_int2002_t(x : std_logic_vector) return int2002_t;
subtype uint2003_t is unsigned(2002 downto 0);
constant uint2003_t_SLV_LEN : integer := 2003;
function uint2003_t_to_slv(x : uint2003_t) return std_logic_vector;
function slv_to_uint2003_t(x : std_logic_vector) return uint2003_t;
subtype int2003_t is signed(2002 downto 0);
constant int2003_t_SLV_LEN : integer := 2003;
function int2003_t_to_slv(x : int2003_t) return std_logic_vector;
function slv_to_int2003_t(x : std_logic_vector) return int2003_t;
subtype uint2004_t is unsigned(2003 downto 0);
constant uint2004_t_SLV_LEN : integer := 2004;
function uint2004_t_to_slv(x : uint2004_t) return std_logic_vector;
function slv_to_uint2004_t(x : std_logic_vector) return uint2004_t;
subtype int2004_t is signed(2003 downto 0);
constant int2004_t_SLV_LEN : integer := 2004;
function int2004_t_to_slv(x : int2004_t) return std_logic_vector;
function slv_to_int2004_t(x : std_logic_vector) return int2004_t;
subtype uint2005_t is unsigned(2004 downto 0);
constant uint2005_t_SLV_LEN : integer := 2005;
function uint2005_t_to_slv(x : uint2005_t) return std_logic_vector;
function slv_to_uint2005_t(x : std_logic_vector) return uint2005_t;
subtype int2005_t is signed(2004 downto 0);
constant int2005_t_SLV_LEN : integer := 2005;
function int2005_t_to_slv(x : int2005_t) return std_logic_vector;
function slv_to_int2005_t(x : std_logic_vector) return int2005_t;
subtype uint2006_t is unsigned(2005 downto 0);
constant uint2006_t_SLV_LEN : integer := 2006;
function uint2006_t_to_slv(x : uint2006_t) return std_logic_vector;
function slv_to_uint2006_t(x : std_logic_vector) return uint2006_t;
subtype int2006_t is signed(2005 downto 0);
constant int2006_t_SLV_LEN : integer := 2006;
function int2006_t_to_slv(x : int2006_t) return std_logic_vector;
function slv_to_int2006_t(x : std_logic_vector) return int2006_t;
subtype uint2007_t is unsigned(2006 downto 0);
constant uint2007_t_SLV_LEN : integer := 2007;
function uint2007_t_to_slv(x : uint2007_t) return std_logic_vector;
function slv_to_uint2007_t(x : std_logic_vector) return uint2007_t;
subtype int2007_t is signed(2006 downto 0);
constant int2007_t_SLV_LEN : integer := 2007;
function int2007_t_to_slv(x : int2007_t) return std_logic_vector;
function slv_to_int2007_t(x : std_logic_vector) return int2007_t;
subtype uint2008_t is unsigned(2007 downto 0);
constant uint2008_t_SLV_LEN : integer := 2008;
function uint2008_t_to_slv(x : uint2008_t) return std_logic_vector;
function slv_to_uint2008_t(x : std_logic_vector) return uint2008_t;
subtype int2008_t is signed(2007 downto 0);
constant int2008_t_SLV_LEN : integer := 2008;
function int2008_t_to_slv(x : int2008_t) return std_logic_vector;
function slv_to_int2008_t(x : std_logic_vector) return int2008_t;
subtype uint2009_t is unsigned(2008 downto 0);
constant uint2009_t_SLV_LEN : integer := 2009;
function uint2009_t_to_slv(x : uint2009_t) return std_logic_vector;
function slv_to_uint2009_t(x : std_logic_vector) return uint2009_t;
subtype int2009_t is signed(2008 downto 0);
constant int2009_t_SLV_LEN : integer := 2009;
function int2009_t_to_slv(x : int2009_t) return std_logic_vector;
function slv_to_int2009_t(x : std_logic_vector) return int2009_t;
subtype uint2010_t is unsigned(2009 downto 0);
constant uint2010_t_SLV_LEN : integer := 2010;
function uint2010_t_to_slv(x : uint2010_t) return std_logic_vector;
function slv_to_uint2010_t(x : std_logic_vector) return uint2010_t;
subtype int2010_t is signed(2009 downto 0);
constant int2010_t_SLV_LEN : integer := 2010;
function int2010_t_to_slv(x : int2010_t) return std_logic_vector;
function slv_to_int2010_t(x : std_logic_vector) return int2010_t;
subtype uint2011_t is unsigned(2010 downto 0);
constant uint2011_t_SLV_LEN : integer := 2011;
function uint2011_t_to_slv(x : uint2011_t) return std_logic_vector;
function slv_to_uint2011_t(x : std_logic_vector) return uint2011_t;
subtype int2011_t is signed(2010 downto 0);
constant int2011_t_SLV_LEN : integer := 2011;
function int2011_t_to_slv(x : int2011_t) return std_logic_vector;
function slv_to_int2011_t(x : std_logic_vector) return int2011_t;
subtype uint2012_t is unsigned(2011 downto 0);
constant uint2012_t_SLV_LEN : integer := 2012;
function uint2012_t_to_slv(x : uint2012_t) return std_logic_vector;
function slv_to_uint2012_t(x : std_logic_vector) return uint2012_t;
subtype int2012_t is signed(2011 downto 0);
constant int2012_t_SLV_LEN : integer := 2012;
function int2012_t_to_slv(x : int2012_t) return std_logic_vector;
function slv_to_int2012_t(x : std_logic_vector) return int2012_t;
subtype uint2013_t is unsigned(2012 downto 0);
constant uint2013_t_SLV_LEN : integer := 2013;
function uint2013_t_to_slv(x : uint2013_t) return std_logic_vector;
function slv_to_uint2013_t(x : std_logic_vector) return uint2013_t;
subtype int2013_t is signed(2012 downto 0);
constant int2013_t_SLV_LEN : integer := 2013;
function int2013_t_to_slv(x : int2013_t) return std_logic_vector;
function slv_to_int2013_t(x : std_logic_vector) return int2013_t;
subtype uint2014_t is unsigned(2013 downto 0);
constant uint2014_t_SLV_LEN : integer := 2014;
function uint2014_t_to_slv(x : uint2014_t) return std_logic_vector;
function slv_to_uint2014_t(x : std_logic_vector) return uint2014_t;
subtype int2014_t is signed(2013 downto 0);
constant int2014_t_SLV_LEN : integer := 2014;
function int2014_t_to_slv(x : int2014_t) return std_logic_vector;
function slv_to_int2014_t(x : std_logic_vector) return int2014_t;
subtype uint2015_t is unsigned(2014 downto 0);
constant uint2015_t_SLV_LEN : integer := 2015;
function uint2015_t_to_slv(x : uint2015_t) return std_logic_vector;
function slv_to_uint2015_t(x : std_logic_vector) return uint2015_t;
subtype int2015_t is signed(2014 downto 0);
constant int2015_t_SLV_LEN : integer := 2015;
function int2015_t_to_slv(x : int2015_t) return std_logic_vector;
function slv_to_int2015_t(x : std_logic_vector) return int2015_t;
subtype uint2016_t is unsigned(2015 downto 0);
constant uint2016_t_SLV_LEN : integer := 2016;
function uint2016_t_to_slv(x : uint2016_t) return std_logic_vector;
function slv_to_uint2016_t(x : std_logic_vector) return uint2016_t;
subtype int2016_t is signed(2015 downto 0);
constant int2016_t_SLV_LEN : integer := 2016;
function int2016_t_to_slv(x : int2016_t) return std_logic_vector;
function slv_to_int2016_t(x : std_logic_vector) return int2016_t;
subtype uint2017_t is unsigned(2016 downto 0);
constant uint2017_t_SLV_LEN : integer := 2017;
function uint2017_t_to_slv(x : uint2017_t) return std_logic_vector;
function slv_to_uint2017_t(x : std_logic_vector) return uint2017_t;
subtype int2017_t is signed(2016 downto 0);
constant int2017_t_SLV_LEN : integer := 2017;
function int2017_t_to_slv(x : int2017_t) return std_logic_vector;
function slv_to_int2017_t(x : std_logic_vector) return int2017_t;
subtype uint2018_t is unsigned(2017 downto 0);
constant uint2018_t_SLV_LEN : integer := 2018;
function uint2018_t_to_slv(x : uint2018_t) return std_logic_vector;
function slv_to_uint2018_t(x : std_logic_vector) return uint2018_t;
subtype int2018_t is signed(2017 downto 0);
constant int2018_t_SLV_LEN : integer := 2018;
function int2018_t_to_slv(x : int2018_t) return std_logic_vector;
function slv_to_int2018_t(x : std_logic_vector) return int2018_t;
subtype uint2019_t is unsigned(2018 downto 0);
constant uint2019_t_SLV_LEN : integer := 2019;
function uint2019_t_to_slv(x : uint2019_t) return std_logic_vector;
function slv_to_uint2019_t(x : std_logic_vector) return uint2019_t;
subtype int2019_t is signed(2018 downto 0);
constant int2019_t_SLV_LEN : integer := 2019;
function int2019_t_to_slv(x : int2019_t) return std_logic_vector;
function slv_to_int2019_t(x : std_logic_vector) return int2019_t;
subtype uint2020_t is unsigned(2019 downto 0);
constant uint2020_t_SLV_LEN : integer := 2020;
function uint2020_t_to_slv(x : uint2020_t) return std_logic_vector;
function slv_to_uint2020_t(x : std_logic_vector) return uint2020_t;
subtype int2020_t is signed(2019 downto 0);
constant int2020_t_SLV_LEN : integer := 2020;
function int2020_t_to_slv(x : int2020_t) return std_logic_vector;
function slv_to_int2020_t(x : std_logic_vector) return int2020_t;
subtype uint2021_t is unsigned(2020 downto 0);
constant uint2021_t_SLV_LEN : integer := 2021;
function uint2021_t_to_slv(x : uint2021_t) return std_logic_vector;
function slv_to_uint2021_t(x : std_logic_vector) return uint2021_t;
subtype int2021_t is signed(2020 downto 0);
constant int2021_t_SLV_LEN : integer := 2021;
function int2021_t_to_slv(x : int2021_t) return std_logic_vector;
function slv_to_int2021_t(x : std_logic_vector) return int2021_t;
subtype uint2022_t is unsigned(2021 downto 0);
constant uint2022_t_SLV_LEN : integer := 2022;
function uint2022_t_to_slv(x : uint2022_t) return std_logic_vector;
function slv_to_uint2022_t(x : std_logic_vector) return uint2022_t;
subtype int2022_t is signed(2021 downto 0);
constant int2022_t_SLV_LEN : integer := 2022;
function int2022_t_to_slv(x : int2022_t) return std_logic_vector;
function slv_to_int2022_t(x : std_logic_vector) return int2022_t;
subtype uint2023_t is unsigned(2022 downto 0);
constant uint2023_t_SLV_LEN : integer := 2023;
function uint2023_t_to_slv(x : uint2023_t) return std_logic_vector;
function slv_to_uint2023_t(x : std_logic_vector) return uint2023_t;
subtype int2023_t is signed(2022 downto 0);
constant int2023_t_SLV_LEN : integer := 2023;
function int2023_t_to_slv(x : int2023_t) return std_logic_vector;
function slv_to_int2023_t(x : std_logic_vector) return int2023_t;
subtype uint2024_t is unsigned(2023 downto 0);
constant uint2024_t_SLV_LEN : integer := 2024;
function uint2024_t_to_slv(x : uint2024_t) return std_logic_vector;
function slv_to_uint2024_t(x : std_logic_vector) return uint2024_t;
subtype int2024_t is signed(2023 downto 0);
constant int2024_t_SLV_LEN : integer := 2024;
function int2024_t_to_slv(x : int2024_t) return std_logic_vector;
function slv_to_int2024_t(x : std_logic_vector) return int2024_t;
subtype uint2025_t is unsigned(2024 downto 0);
constant uint2025_t_SLV_LEN : integer := 2025;
function uint2025_t_to_slv(x : uint2025_t) return std_logic_vector;
function slv_to_uint2025_t(x : std_logic_vector) return uint2025_t;
subtype int2025_t is signed(2024 downto 0);
constant int2025_t_SLV_LEN : integer := 2025;
function int2025_t_to_slv(x : int2025_t) return std_logic_vector;
function slv_to_int2025_t(x : std_logic_vector) return int2025_t;
subtype uint2026_t is unsigned(2025 downto 0);
constant uint2026_t_SLV_LEN : integer := 2026;
function uint2026_t_to_slv(x : uint2026_t) return std_logic_vector;
function slv_to_uint2026_t(x : std_logic_vector) return uint2026_t;
subtype int2026_t is signed(2025 downto 0);
constant int2026_t_SLV_LEN : integer := 2026;
function int2026_t_to_slv(x : int2026_t) return std_logic_vector;
function slv_to_int2026_t(x : std_logic_vector) return int2026_t;
subtype uint2027_t is unsigned(2026 downto 0);
constant uint2027_t_SLV_LEN : integer := 2027;
function uint2027_t_to_slv(x : uint2027_t) return std_logic_vector;
function slv_to_uint2027_t(x : std_logic_vector) return uint2027_t;
subtype int2027_t is signed(2026 downto 0);
constant int2027_t_SLV_LEN : integer := 2027;
function int2027_t_to_slv(x : int2027_t) return std_logic_vector;
function slv_to_int2027_t(x : std_logic_vector) return int2027_t;
subtype uint2028_t is unsigned(2027 downto 0);
constant uint2028_t_SLV_LEN : integer := 2028;
function uint2028_t_to_slv(x : uint2028_t) return std_logic_vector;
function slv_to_uint2028_t(x : std_logic_vector) return uint2028_t;
subtype int2028_t is signed(2027 downto 0);
constant int2028_t_SLV_LEN : integer := 2028;
function int2028_t_to_slv(x : int2028_t) return std_logic_vector;
function slv_to_int2028_t(x : std_logic_vector) return int2028_t;
subtype uint2029_t is unsigned(2028 downto 0);
constant uint2029_t_SLV_LEN : integer := 2029;
function uint2029_t_to_slv(x : uint2029_t) return std_logic_vector;
function slv_to_uint2029_t(x : std_logic_vector) return uint2029_t;
subtype int2029_t is signed(2028 downto 0);
constant int2029_t_SLV_LEN : integer := 2029;
function int2029_t_to_slv(x : int2029_t) return std_logic_vector;
function slv_to_int2029_t(x : std_logic_vector) return int2029_t;
subtype uint2030_t is unsigned(2029 downto 0);
constant uint2030_t_SLV_LEN : integer := 2030;
function uint2030_t_to_slv(x : uint2030_t) return std_logic_vector;
function slv_to_uint2030_t(x : std_logic_vector) return uint2030_t;
subtype int2030_t is signed(2029 downto 0);
constant int2030_t_SLV_LEN : integer := 2030;
function int2030_t_to_slv(x : int2030_t) return std_logic_vector;
function slv_to_int2030_t(x : std_logic_vector) return int2030_t;
subtype uint2031_t is unsigned(2030 downto 0);
constant uint2031_t_SLV_LEN : integer := 2031;
function uint2031_t_to_slv(x : uint2031_t) return std_logic_vector;
function slv_to_uint2031_t(x : std_logic_vector) return uint2031_t;
subtype int2031_t is signed(2030 downto 0);
constant int2031_t_SLV_LEN : integer := 2031;
function int2031_t_to_slv(x : int2031_t) return std_logic_vector;
function slv_to_int2031_t(x : std_logic_vector) return int2031_t;
subtype uint2032_t is unsigned(2031 downto 0);
constant uint2032_t_SLV_LEN : integer := 2032;
function uint2032_t_to_slv(x : uint2032_t) return std_logic_vector;
function slv_to_uint2032_t(x : std_logic_vector) return uint2032_t;
subtype int2032_t is signed(2031 downto 0);
constant int2032_t_SLV_LEN : integer := 2032;
function int2032_t_to_slv(x : int2032_t) return std_logic_vector;
function slv_to_int2032_t(x : std_logic_vector) return int2032_t;
subtype uint2033_t is unsigned(2032 downto 0);
constant uint2033_t_SLV_LEN : integer := 2033;
function uint2033_t_to_slv(x : uint2033_t) return std_logic_vector;
function slv_to_uint2033_t(x : std_logic_vector) return uint2033_t;
subtype int2033_t is signed(2032 downto 0);
constant int2033_t_SLV_LEN : integer := 2033;
function int2033_t_to_slv(x : int2033_t) return std_logic_vector;
function slv_to_int2033_t(x : std_logic_vector) return int2033_t;
subtype uint2034_t is unsigned(2033 downto 0);
constant uint2034_t_SLV_LEN : integer := 2034;
function uint2034_t_to_slv(x : uint2034_t) return std_logic_vector;
function slv_to_uint2034_t(x : std_logic_vector) return uint2034_t;
subtype int2034_t is signed(2033 downto 0);
constant int2034_t_SLV_LEN : integer := 2034;
function int2034_t_to_slv(x : int2034_t) return std_logic_vector;
function slv_to_int2034_t(x : std_logic_vector) return int2034_t;
subtype uint2035_t is unsigned(2034 downto 0);
constant uint2035_t_SLV_LEN : integer := 2035;
function uint2035_t_to_slv(x : uint2035_t) return std_logic_vector;
function slv_to_uint2035_t(x : std_logic_vector) return uint2035_t;
subtype int2035_t is signed(2034 downto 0);
constant int2035_t_SLV_LEN : integer := 2035;
function int2035_t_to_slv(x : int2035_t) return std_logic_vector;
function slv_to_int2035_t(x : std_logic_vector) return int2035_t;
subtype uint2036_t is unsigned(2035 downto 0);
constant uint2036_t_SLV_LEN : integer := 2036;
function uint2036_t_to_slv(x : uint2036_t) return std_logic_vector;
function slv_to_uint2036_t(x : std_logic_vector) return uint2036_t;
subtype int2036_t is signed(2035 downto 0);
constant int2036_t_SLV_LEN : integer := 2036;
function int2036_t_to_slv(x : int2036_t) return std_logic_vector;
function slv_to_int2036_t(x : std_logic_vector) return int2036_t;
subtype uint2037_t is unsigned(2036 downto 0);
constant uint2037_t_SLV_LEN : integer := 2037;
function uint2037_t_to_slv(x : uint2037_t) return std_logic_vector;
function slv_to_uint2037_t(x : std_logic_vector) return uint2037_t;
subtype int2037_t is signed(2036 downto 0);
constant int2037_t_SLV_LEN : integer := 2037;
function int2037_t_to_slv(x : int2037_t) return std_logic_vector;
function slv_to_int2037_t(x : std_logic_vector) return int2037_t;
subtype uint2038_t is unsigned(2037 downto 0);
constant uint2038_t_SLV_LEN : integer := 2038;
function uint2038_t_to_slv(x : uint2038_t) return std_logic_vector;
function slv_to_uint2038_t(x : std_logic_vector) return uint2038_t;
subtype int2038_t is signed(2037 downto 0);
constant int2038_t_SLV_LEN : integer := 2038;
function int2038_t_to_slv(x : int2038_t) return std_logic_vector;
function slv_to_int2038_t(x : std_logic_vector) return int2038_t;
subtype uint2039_t is unsigned(2038 downto 0);
constant uint2039_t_SLV_LEN : integer := 2039;
function uint2039_t_to_slv(x : uint2039_t) return std_logic_vector;
function slv_to_uint2039_t(x : std_logic_vector) return uint2039_t;
subtype int2039_t is signed(2038 downto 0);
constant int2039_t_SLV_LEN : integer := 2039;
function int2039_t_to_slv(x : int2039_t) return std_logic_vector;
function slv_to_int2039_t(x : std_logic_vector) return int2039_t;
subtype uint2040_t is unsigned(2039 downto 0);
constant uint2040_t_SLV_LEN : integer := 2040;
function uint2040_t_to_slv(x : uint2040_t) return std_logic_vector;
function slv_to_uint2040_t(x : std_logic_vector) return uint2040_t;
subtype int2040_t is signed(2039 downto 0);
constant int2040_t_SLV_LEN : integer := 2040;
function int2040_t_to_slv(x : int2040_t) return std_logic_vector;
function slv_to_int2040_t(x : std_logic_vector) return int2040_t;
subtype uint2041_t is unsigned(2040 downto 0);
constant uint2041_t_SLV_LEN : integer := 2041;
function uint2041_t_to_slv(x : uint2041_t) return std_logic_vector;
function slv_to_uint2041_t(x : std_logic_vector) return uint2041_t;
subtype int2041_t is signed(2040 downto 0);
constant int2041_t_SLV_LEN : integer := 2041;
function int2041_t_to_slv(x : int2041_t) return std_logic_vector;
function slv_to_int2041_t(x : std_logic_vector) return int2041_t;
subtype uint2042_t is unsigned(2041 downto 0);
constant uint2042_t_SLV_LEN : integer := 2042;
function uint2042_t_to_slv(x : uint2042_t) return std_logic_vector;
function slv_to_uint2042_t(x : std_logic_vector) return uint2042_t;
subtype int2042_t is signed(2041 downto 0);
constant int2042_t_SLV_LEN : integer := 2042;
function int2042_t_to_slv(x : int2042_t) return std_logic_vector;
function slv_to_int2042_t(x : std_logic_vector) return int2042_t;
subtype uint2043_t is unsigned(2042 downto 0);
constant uint2043_t_SLV_LEN : integer := 2043;
function uint2043_t_to_slv(x : uint2043_t) return std_logic_vector;
function slv_to_uint2043_t(x : std_logic_vector) return uint2043_t;
subtype int2043_t is signed(2042 downto 0);
constant int2043_t_SLV_LEN : integer := 2043;
function int2043_t_to_slv(x : int2043_t) return std_logic_vector;
function slv_to_int2043_t(x : std_logic_vector) return int2043_t;
subtype uint2044_t is unsigned(2043 downto 0);
constant uint2044_t_SLV_LEN : integer := 2044;
function uint2044_t_to_slv(x : uint2044_t) return std_logic_vector;
function slv_to_uint2044_t(x : std_logic_vector) return uint2044_t;
subtype int2044_t is signed(2043 downto 0);
constant int2044_t_SLV_LEN : integer := 2044;
function int2044_t_to_slv(x : int2044_t) return std_logic_vector;
function slv_to_int2044_t(x : std_logic_vector) return int2044_t;
subtype uint2045_t is unsigned(2044 downto 0);
constant uint2045_t_SLV_LEN : integer := 2045;
function uint2045_t_to_slv(x : uint2045_t) return std_logic_vector;
function slv_to_uint2045_t(x : std_logic_vector) return uint2045_t;
subtype int2045_t is signed(2044 downto 0);
constant int2045_t_SLV_LEN : integer := 2045;
function int2045_t_to_slv(x : int2045_t) return std_logic_vector;
function slv_to_int2045_t(x : std_logic_vector) return int2045_t;
subtype uint2046_t is unsigned(2045 downto 0);
constant uint2046_t_SLV_LEN : integer := 2046;
function uint2046_t_to_slv(x : uint2046_t) return std_logic_vector;
function slv_to_uint2046_t(x : std_logic_vector) return uint2046_t;
subtype int2046_t is signed(2045 downto 0);
constant int2046_t_SLV_LEN : integer := 2046;
function int2046_t_to_slv(x : int2046_t) return std_logic_vector;
function slv_to_int2046_t(x : std_logic_vector) return int2046_t;
subtype uint2047_t is unsigned(2046 downto 0);
constant uint2047_t_SLV_LEN : integer := 2047;
function uint2047_t_to_slv(x : uint2047_t) return std_logic_vector;
function slv_to_uint2047_t(x : std_logic_vector) return uint2047_t;
subtype int2047_t is signed(2046 downto 0);
constant int2047_t_SLV_LEN : integer := 2047;
function int2047_t_to_slv(x : int2047_t) return std_logic_vector;
function slv_to_int2047_t(x : std_logic_vector) return int2047_t;
subtype uint2048_t is unsigned(2047 downto 0);
constant uint2048_t_SLV_LEN : integer := 2048;
function uint2048_t_to_slv(x : uint2048_t) return std_logic_vector;
function slv_to_uint2048_t(x : std_logic_vector) return uint2048_t;
subtype int2048_t is signed(2047 downto 0);
constant int2048_t_SLV_LEN : integer := 2048;
function int2048_t_to_slv(x : int2048_t) return std_logic_vector;
function slv_to_int2048_t(x : std_logic_vector) return int2048_t;

  type byte_array_t is array (natural range <>) of unsigned(7 downto 0);
  function to_byte_array(s : string; constant len : natural) return byte_array_t;
  
  function resize_float_e_m_t(
    x : std_logic_vector; 
    in_exponent_width : integer;
    in_mantissa_width : integer;
    out_exponent_width : integer;
    out_mantissa_width : integer) return std_logic_vector; 
   
  type chacha20_decrypt_state_t is (
    
      POLY_KEY,
      PLAINTEXT
  );
  
function chacha20_decrypt_state_t_to_slv(e : chacha20_decrypt_state_t) return std_logic_vector;

  type prep_auth_data_state_t is (
    
      IDLE,
      AAD,
      CIPHERTEXT,
      LENGTHS
  );
  
function prep_auth_data_state_t_to_slv(e : prep_auth_data_state_t) return std_logic_vector;

  type poly1305_state_t is (
    
      IDLE,
      START_ITER,
      FINISH_ITER,
      A_PLUS_S,
      OUTPUT_AUTH_TAG
  );
  
function poly1305_state_t_to_slv(e : poly1305_state_t) return std_logic_vector;

  type poly1305_verify_state_t is (
    
      TAKE_AUTH_TAG,
      TAKE_CALC_TAG,
      COMPARE_TAGS,
      OUTPUT_COMPARE_RESULT
  );
  
function poly1305_verify_state_t_to_slv(e : poly1305_verify_state_t) return std_logic_vector;

  type strip_auth_tag_state_t is (
    
      CIPHERTEXT_PASS,
      AUTH_TAG_EXTRACTION
  );
  
function strip_auth_tag_state_t_to_slv(e : strip_auth_tag_state_t) return std_logic_vector;

  type wait_to_verify_state_t is (
    
      WAIT_TO_VERIFY_BIT,
      OUTPUT_PLAINTEXT
  );
  
function wait_to_verify_state_t_to_slv(e : wait_to_verify_state_t) return std_logic_vector;
subtype uint8_t_16 is byte_array_t(0 to 15);
constant uint8_t_16_SLV_LEN : integer := 8 * 16;

      function uint8_t_16_to_slv(data : uint8_t_16) return std_logic_vector;

      function slv_to_uint8_t_16(data : std_logic_vector) return uint8_t_16;
type uint64_t_5 is array(0 to 4) of unsigned(63 downto 0);
constant uint64_t_5_SLV_LEN : integer := 64 * 5;

      function uint64_t_5_to_slv(data : uint64_t_5) return std_logic_vector;

      function slv_to_uint64_t_5(data : std_logic_vector) return uint64_t_5;
subtype uint8_t_32 is byte_array_t(0 to 31);
constant uint8_t_32_SLV_LEN : integer := 8 * 32;

      function uint8_t_32_to_slv(data : uint8_t_32) return std_logic_vector;

      function slv_to_uint8_t_32(data : std_logic_vector) return uint8_t_32;
subtype uint8_t_12 is byte_array_t(0 to 11);
constant uint8_t_12_SLV_LEN : integer := 8 * 12;

      function uint8_t_12_to_slv(data : uint8_t_12) return std_logic_vector;

      function slv_to_uint8_t_12(data : std_logic_vector) return uint8_t_12;
type uint1_t_64 is array(0 to 63) of unsigned(0 downto 0);
constant uint1_t_64_SLV_LEN : integer := 1 * 64;

      function uint1_t_64_to_slv(data : uint1_t_64) return std_logic_vector;

      function slv_to_uint1_t_64(data : std_logic_vector) return uint1_t_64;
type uint1_t_16 is array(0 to 15) of unsigned(0 downto 0);
constant uint1_t_16_SLV_LEN : integer := 1 * 16;

      function uint1_t_16_to_slv(data : uint1_t_16) return std_logic_vector;

      function slv_to_uint1_t_16(data : std_logic_vector) return uint1_t_16;
type uint32_t_8 is array(0 to 7) of unsigned(31 downto 0);
constant uint32_t_8_SLV_LEN : integer := 32 * 8;

      function uint32_t_8_to_slv(data : uint32_t_8) return std_logic_vector;

      function slv_to_uint32_t_8(data : std_logic_vector) return uint32_t_8;
type uint32_t_3 is array(0 to 2) of unsigned(31 downto 0);
constant uint32_t_3_SLV_LEN : integer := 32 * 3;

      function uint32_t_3_to_slv(data : uint32_t_3) return std_logic_vector;

      function slv_to_uint32_t_3(data : std_logic_vector) return uint32_t_3;
subtype uint8_t_64 is byte_array_t(0 to 63);
constant uint8_t_64_SLV_LEN : integer := 8 * 64;

      function uint8_t_64_to_slv(data : uint8_t_64) return std_logic_vector;

      function slv_to_uint8_t_64(data : std_logic_vector) return uint8_t_64;
subtype uint8_t_8 is byte_array_t(0 to 7);
constant uint8_t_8_SLV_LEN : integer := 8 * 8;

      function uint8_t_8_to_slv(data : uint8_t_8) return std_logic_vector;

      function slv_to_uint8_t_8(data : std_logic_vector) return uint8_t_8;
subtype uint8_t_40 is byte_array_t(0 to 39);
constant uint8_t_40_SLV_LEN : integer := 8 * 40;

      function uint8_t_40_to_slv(data : uint8_t_40) return std_logic_vector;

      function slv_to_uint8_t_40(data : std_logic_vector) return uint8_t_40;
subtype char_128 is byte_array_t(0 to 127);
constant char_128_SLV_LEN : integer := 8 * 128;

      function char_128_to_slv(data : char_128) return std_logic_vector;

      function slv_to_char_128(data : std_logic_vector) return char_128;
type char_2_128 is array(0 to 1) of char_128;
constant char_2_128_SLV_LEN : integer := char_128_SLV_LEN * 2;

      function char_2_128_to_slv(data : char_2_128) return std_logic_vector;

      function slv_to_char_2_128(data : std_logic_vector) return char_2_128;
type uint32_t_2 is array(0 to 1) of unsigned(31 downto 0);
constant uint32_t_2_SLV_LEN : integer := 32 * 2;

      function uint32_t_2_to_slv(data : uint32_t_2) return std_logic_vector;

      function slv_to_uint32_t_2(data : std_logic_vector) return uint32_t_2;
subtype uint8_t_144 is byte_array_t(0 to 143);
constant uint8_t_144_SLV_LEN : integer := 8 * 144;

      function uint8_t_144_to_slv(data : uint8_t_144) return std_logic_vector;

      function slv_to_uint8_t_144(data : std_logic_vector) return uint8_t_144;
type uint8_t_2_144 is array(0 to 1) of uint8_t_144;
constant uint8_t_2_144_SLV_LEN : integer := uint8_t_144_SLV_LEN * 2;

      function uint8_t_2_144_to_slv(data : uint8_t_2_144) return std_logic_vector;

      function slv_to_uint8_t_2_144(data : std_logic_vector) return uint8_t_2_144;
subtype uint8_t_1 is byte_array_t(0 to 0);
constant uint8_t_1_SLV_LEN : integer := 8 * 1;

      function uint8_t_1_to_slv(data : uint8_t_1) return std_logic_vector;

      function slv_to_uint8_t_1(data : std_logic_vector) return uint8_t_1;
type uint1_t_1 is array(0 to 0) of unsigned(0 downto 0);
constant uint1_t_1_SLV_LEN : integer := 1 * 1;

      function uint1_t_1_to_slv(data : uint1_t_1) return std_logic_vector;

      function slv_to_uint1_t_1(data : std_logic_vector) return uint1_t_1;
subtype uint8_t_2 is byte_array_t(0 to 1);
constant uint8_t_2_SLV_LEN : integer := 8 * 2;

      function uint8_t_2_to_slv(data : uint8_t_2) return std_logic_vector;

      function slv_to_uint8_t_2(data : std_logic_vector) return uint8_t_2;
type uint1_t_2 is array(0 to 1) of unsigned(0 downto 0);
constant uint1_t_2_SLV_LEN : integer := 1 * 2;

      function uint1_t_2_to_slv(data : uint1_t_2) return std_logic_vector;

      function slv_to_uint1_t_2(data : std_logic_vector) return uint1_t_2;
subtype uint8_t_4 is byte_array_t(0 to 3);
constant uint8_t_4_SLV_LEN : integer := 8 * 4;

      function uint8_t_4_to_slv(data : uint8_t_4) return std_logic_vector;

      function slv_to_uint8_t_4(data : std_logic_vector) return uint8_t_4;
type uint1_t_4 is array(0 to 3) of unsigned(0 downto 0);
constant uint1_t_4_SLV_LEN : integer := 1 * 4;

      function uint1_t_4_to_slv(data : uint1_t_4) return std_logic_vector;

      function slv_to_uint1_t_4(data : std_logic_vector) return uint1_t_4;
type uint1_t_8 is array(0 to 7) of unsigned(0 downto 0);
constant uint1_t_8_SLV_LEN : integer := 1 * 8;

      function uint1_t_8_to_slv(data : uint1_t_8) return std_logic_vector;

      function slv_to_uint1_t_8(data : std_logic_vector) return uint1_t_8;
type uint1_t_32 is array(0 to 31) of unsigned(0 downto 0);
constant uint1_t_32_SLV_LEN : integer := 1 * 32;

      function uint1_t_32_to_slv(data : uint1_t_32) return std_logic_vector;

      function slv_to_uint1_t_32(data : std_logic_vector) return uint1_t_32;
type uint32_t_16 is array(0 to 15) of unsigned(31 downto 0);
constant uint32_t_16_SLV_LEN : integer := 32 * 16;

      function uint32_t_16_to_slv(data : uint32_t_16) return std_logic_vector;

      function slv_to_uint32_t_16(data : std_logic_vector) return uint32_t_16;

  type axis8_t is record
  
    tdata : uint8_t_1;
    tkeep : uint1_t_1;
    tlast : unsigned(0 downto 0);
  end record;
  
  constant axis8_t_NULL : axis8_t := (
  
    tdata => (others => to_unsigned(0, 8)),
    tkeep => (others => to_unsigned(0, 1)),
    tlast => to_unsigned(0, 1)
  );
  
  constant axis8_t_SLV_LEN : integer := (
  uint8_t_1_SLV_LEN+uint1_t_1_SLV_LEN+1
  );
  
  function axis8_t_to_slv(data : axis8_t) return std_logic_vector;

  function slv_to_axis8_t(data : std_logic_vector) return axis8_t;

  type axis8_t_stream_t is record
  
    data : axis8_t;
    valid : unsigned(0 downto 0);
  end record;
  
  constant axis8_t_stream_t_NULL : axis8_t_stream_t := (
  
    data => axis8_t_NULL,
    valid => to_unsigned(0, 1)
  );
  
  constant axis8_t_stream_t_SLV_LEN : integer := (
  axis8_t_SLV_LEN+1
  );
  
  function axis8_t_stream_t_to_slv(data : axis8_t_stream_t) return std_logic_vector;

  function slv_to_axis8_t_stream_t(data : std_logic_vector) return axis8_t_stream_t;

  type axis16_t is record
  
    tdata : uint8_t_2;
    tkeep : uint1_t_2;
    tlast : unsigned(0 downto 0);
  end record;
  
  constant axis16_t_NULL : axis16_t := (
  
    tdata => (others => to_unsigned(0, 8)),
    tkeep => (others => to_unsigned(0, 1)),
    tlast => to_unsigned(0, 1)
  );
  
  constant axis16_t_SLV_LEN : integer := (
  uint8_t_2_SLV_LEN+uint1_t_2_SLV_LEN+1
  );
  
  function axis16_t_to_slv(data : axis16_t) return std_logic_vector;

  function slv_to_axis16_t(data : std_logic_vector) return axis16_t;

  type axis16_t_stream_t is record
  
    data : axis16_t;
    valid : unsigned(0 downto 0);
  end record;
  
  constant axis16_t_stream_t_NULL : axis16_t_stream_t := (
  
    data => axis16_t_NULL,
    valid => to_unsigned(0, 1)
  );
  
  constant axis16_t_stream_t_SLV_LEN : integer := (
  axis16_t_SLV_LEN+1
  );
  
  function axis16_t_stream_t_to_slv(data : axis16_t_stream_t) return std_logic_vector;

  function slv_to_axis16_t_stream_t(data : std_logic_vector) return axis16_t_stream_t;

  type axis32_t is record
  
    tdata : uint8_t_4;
    tkeep : uint1_t_4;
    tlast : unsigned(0 downto 0);
  end record;
  
  constant axis32_t_NULL : axis32_t := (
  
    tdata => (others => to_unsigned(0, 8)),
    tkeep => (others => to_unsigned(0, 1)),
    tlast => to_unsigned(0, 1)
  );
  
  constant axis32_t_SLV_LEN : integer := (
  uint8_t_4_SLV_LEN+uint1_t_4_SLV_LEN+1
  );
  
  function axis32_t_to_slv(data : axis32_t) return std_logic_vector;

  function slv_to_axis32_t(data : std_logic_vector) return axis32_t;

  type axis32_t_stream_t is record
  
    data : axis32_t;
    valid : unsigned(0 downto 0);
  end record;
  
  constant axis32_t_stream_t_NULL : axis32_t_stream_t := (
  
    data => axis32_t_NULL,
    valid => to_unsigned(0, 1)
  );
  
  constant axis32_t_stream_t_SLV_LEN : integer := (
  axis32_t_SLV_LEN+1
  );
  
  function axis32_t_stream_t_to_slv(data : axis32_t_stream_t) return std_logic_vector;

  function slv_to_axis32_t_stream_t(data : std_logic_vector) return axis32_t_stream_t;

  type axis64_t is record
  
    tdata : uint8_t_8;
    tkeep : uint1_t_8;
    tlast : unsigned(0 downto 0);
  end record;
  
  constant axis64_t_NULL : axis64_t := (
  
    tdata => (others => to_unsigned(0, 8)),
    tkeep => (others => to_unsigned(0, 1)),
    tlast => to_unsigned(0, 1)
  );
  
  constant axis64_t_SLV_LEN : integer := (
  uint8_t_8_SLV_LEN+uint1_t_8_SLV_LEN+1
  );
  
  function axis64_t_to_slv(data : axis64_t) return std_logic_vector;

  function slv_to_axis64_t(data : std_logic_vector) return axis64_t;

  type axis64_t_stream_t is record
  
    data : axis64_t;
    valid : unsigned(0 downto 0);
  end record;
  
  constant axis64_t_stream_t_NULL : axis64_t_stream_t := (
  
    data => axis64_t_NULL,
    valid => to_unsigned(0, 1)
  );
  
  constant axis64_t_stream_t_SLV_LEN : integer := (
  axis64_t_SLV_LEN+1
  );
  
  function axis64_t_stream_t_to_slv(data : axis64_t_stream_t) return std_logic_vector;

  function slv_to_axis64_t_stream_t(data : std_logic_vector) return axis64_t_stream_t;

  type axis128_t is record
  
    tdata : uint8_t_16;
    tkeep : uint1_t_16;
    tlast : unsigned(0 downto 0);
  end record;
  
  constant axis128_t_NULL : axis128_t := (
  
    tdata => (others => to_unsigned(0, 8)),
    tkeep => (others => to_unsigned(0, 1)),
    tlast => to_unsigned(0, 1)
  );
  
  constant axis128_t_SLV_LEN : integer := (
  uint8_t_16_SLV_LEN+uint1_t_16_SLV_LEN+1
  );
  
  function axis128_t_to_slv(data : axis128_t) return std_logic_vector;

  function slv_to_axis128_t(data : std_logic_vector) return axis128_t;

  type axis128_t_stream_t is record
  
    data : axis128_t;
    valid : unsigned(0 downto 0);
  end record;
  
  constant axis128_t_stream_t_NULL : axis128_t_stream_t := (
  
    data => axis128_t_NULL,
    valid => to_unsigned(0, 1)
  );
  
  constant axis128_t_stream_t_SLV_LEN : integer := (
  axis128_t_SLV_LEN+1
  );
  
  function axis128_t_stream_t_to_slv(data : axis128_t_stream_t) return std_logic_vector;

  function slv_to_axis128_t_stream_t(data : std_logic_vector) return axis128_t_stream_t;

  type axis256_t is record
  
    tdata : uint8_t_32;
    tkeep : uint1_t_32;
    tlast : unsigned(0 downto 0);
  end record;
  
  constant axis256_t_NULL : axis256_t := (
  
    tdata => (others => to_unsigned(0, 8)),
    tkeep => (others => to_unsigned(0, 1)),
    tlast => to_unsigned(0, 1)
  );
  
  constant axis256_t_SLV_LEN : integer := (
  uint8_t_32_SLV_LEN+uint1_t_32_SLV_LEN+1
  );
  
  function axis256_t_to_slv(data : axis256_t) return std_logic_vector;

  function slv_to_axis256_t(data : std_logic_vector) return axis256_t;

  type axis256_t_stream_t is record
  
    data : axis256_t;
    valid : unsigned(0 downto 0);
  end record;
  
  constant axis256_t_stream_t_NULL : axis256_t_stream_t := (
  
    data => axis256_t_NULL,
    valid => to_unsigned(0, 1)
  );
  
  constant axis256_t_stream_t_SLV_LEN : integer := (
  axis256_t_SLV_LEN+1
  );
  
  function axis256_t_stream_t_to_slv(data : axis256_t_stream_t) return std_logic_vector;

  function slv_to_axis256_t_stream_t(data : std_logic_vector) return axis256_t_stream_t;

  type axis512_t is record
  
    tdata : uint8_t_64;
    tkeep : uint1_t_64;
    tlast : unsigned(0 downto 0);
  end record;
  
  constant axis512_t_NULL : axis512_t := (
  
    tdata => (others => to_unsigned(0, 8)),
    tkeep => (others => to_unsigned(0, 1)),
    tlast => to_unsigned(0, 1)
  );
  
  constant axis512_t_SLV_LEN : integer := (
  uint8_t_64_SLV_LEN+uint1_t_64_SLV_LEN+1
  );
  
  function axis512_t_to_slv(data : axis512_t) return std_logic_vector;

  function slv_to_axis512_t(data : std_logic_vector) return axis512_t;

  type axis512_t_stream_t is record
  
    data : axis512_t;
    valid : unsigned(0 downto 0);
  end record;
  
  constant axis512_t_stream_t_NULL : axis512_t_stream_t := (
  
    data => axis512_t_NULL,
    valid => to_unsigned(0, 1)
  );
  
  constant axis512_t_stream_t_SLV_LEN : integer := (
  axis512_t_SLV_LEN+1
  );
  
  function axis512_t_stream_t_to_slv(data : axis512_t_stream_t) return std_logic_vector;

  function slv_to_axis512_t_stream_t(data : std_logic_vector) return axis512_t_stream_t;

  type axis8_to_axis32_t is record
  
    axis_out : axis32_t_stream_t;
    axis_in_ready : unsigned(0 downto 0);
  end record;
  
  constant axis8_to_axis32_t_NULL : axis8_to_axis32_t := (
  
    axis_out => axis32_t_stream_t_NULL,
    axis_in_ready => to_unsigned(0, 1)
  );
  
  constant axis8_to_axis32_t_SLV_LEN : integer := (
  axis32_t_stream_t_SLV_LEN+1
  );
  
  function axis8_to_axis32_t_to_slv(data : axis8_to_axis32_t) return std_logic_vector;

  function slv_to_axis8_to_axis32_t(data : std_logic_vector) return axis8_to_axis32_t;

  type axis32_to_axis8_t is record
  
    axis_out : axis8_t_stream_t;
    axis_in_ready : unsigned(0 downto 0);
  end record;
  
  constant axis32_to_axis8_t_NULL : axis32_to_axis8_t := (
  
    axis_out => axis8_t_stream_t_NULL,
    axis_in_ready => to_unsigned(0, 1)
  );
  
  constant axis32_to_axis8_t_SLV_LEN : integer := (
  axis8_t_stream_t_SLV_LEN+1
  );
  
  function axis32_to_axis8_t_to_slv(data : axis32_to_axis8_t) return std_logic_vector;

  function slv_to_axis32_to_axis8_t(data : std_logic_vector) return axis32_to_axis8_t;

  type axis128_to_axis512_t is record
  
    axis_out : axis512_t_stream_t;
    axis_in_ready : unsigned(0 downto 0);
  end record;
  
  constant axis128_to_axis512_t_NULL : axis128_to_axis512_t := (
  
    axis_out => axis512_t_stream_t_NULL,
    axis_in_ready => to_unsigned(0, 1)
  );
  
  constant axis128_to_axis512_t_SLV_LEN : integer := (
  axis512_t_stream_t_SLV_LEN+1
  );
  
  function axis128_to_axis512_t_to_slv(data : axis128_to_axis512_t) return std_logic_vector;

  function slv_to_axis128_to_axis512_t(data : std_logic_vector) return axis128_to_axis512_t;

  type axis512_to_axis128_t is record
  
    axis_out : axis128_t_stream_t;
    axis_in_ready : unsigned(0 downto 0);
  end record;
  
  constant axis512_to_axis128_t_NULL : axis512_to_axis128_t := (
  
    axis_out => axis128_t_stream_t_NULL,
    axis_in_ready => to_unsigned(0, 1)
  );
  
  constant axis512_to_axis128_t_SLV_LEN : integer := (
  axis128_t_stream_t_SLV_LEN+1
  );
  
  function axis512_to_axis128_t_to_slv(data : axis512_to_axis128_t) return std_logic_vector;

  function slv_to_axis512_to_axis128_t(data : std_logic_vector) return axis512_to_axis128_t;

  type axis8_max_len_limiter_t is record
  
    out_stream : axis8_t_stream_t;
    ready_for_in_stream : unsigned(0 downto 0);
  end record;
  
  constant axis8_max_len_limiter_t_NULL : axis8_max_len_limiter_t := (
  
    out_stream => axis8_t_stream_t_NULL,
    ready_for_in_stream => to_unsigned(0, 1)
  );
  
  constant axis8_max_len_limiter_t_SLV_LEN : integer := (
  axis8_t_stream_t_SLV_LEN+1
  );
  
  function axis8_max_len_limiter_t_to_slv(data : axis8_max_len_limiter_t) return std_logic_vector;

  function slv_to_axis8_max_len_limiter_t(data : std_logic_vector) return axis8_max_len_limiter_t;

  type axis32_max_len_limiter_t is record
  
    out_stream : axis32_t_stream_t;
    ready_for_in_stream : unsigned(0 downto 0);
  end record;
  
  constant axis32_max_len_limiter_t_NULL : axis32_max_len_limiter_t := (
  
    out_stream => axis32_t_stream_t_NULL,
    ready_for_in_stream => to_unsigned(0, 1)
  );
  
  constant axis32_max_len_limiter_t_SLV_LEN : integer := (
  axis32_t_stream_t_SLV_LEN+1
  );
  
  function axis32_max_len_limiter_t_to_slv(data : axis32_max_len_limiter_t) return std_logic_vector;

  function slv_to_axis32_max_len_limiter_t(data : std_logic_vector) return axis32_max_len_limiter_t;

  type chacha20_state is record
  
    state : uint32_t_16;
  end record;
  
  constant chacha20_state_NULL : chacha20_state := (
  
    state => (others => to_unsigned(0, 32))
  );
  
  constant chacha20_state_SLV_LEN : integer := (
  uint32_t_16_SLV_LEN
  );
  
  function chacha20_state_to_slv(data : chacha20_state) return std_logic_vector;

  function slv_to_chacha20_state(data : std_logic_vector) return chacha20_state;

  type chacha20_decrypt_loop_body_in_t is record
  
    axis_in : axis512_t;
    key : uint8_t_32;
    nonce : uint8_t_12;
    counter : unsigned(31 downto 0);
  end record;
  
  constant chacha20_decrypt_loop_body_in_t_NULL : chacha20_decrypt_loop_body_in_t := (
  
    axis_in => axis512_t_NULL,
    key => (others => to_unsigned(0, 8)),
    nonce => (others => to_unsigned(0, 8)),
    counter => to_unsigned(0, 32)
  );
  
  constant chacha20_decrypt_loop_body_in_t_SLV_LEN : integer := (
  axis512_t_SLV_LEN+uint8_t_32_SLV_LEN+uint8_t_12_SLV_LEN+32
  );
  
  function chacha20_decrypt_loop_body_in_t_to_slv(data : chacha20_decrypt_loop_body_in_t) return std_logic_vector;

  function slv_to_chacha20_decrypt_loop_body_in_t(data : std_logic_vector) return chacha20_decrypt_loop_body_in_t;

  type chacha20_decrypt_loop_body_in_t_stream_t is record
  
    data : chacha20_decrypt_loop_body_in_t;
    valid : unsigned(0 downto 0);
  end record;
  
  constant chacha20_decrypt_loop_body_in_t_stream_t_NULL : chacha20_decrypt_loop_body_in_t_stream_t := (
  
    data => chacha20_decrypt_loop_body_in_t_NULL,
    valid => to_unsigned(0, 1)
  );
  
  constant chacha20_decrypt_loop_body_in_t_stream_t_SLV_LEN : integer := (
  chacha20_decrypt_loop_body_in_t_SLV_LEN+1
  );
  
  function chacha20_decrypt_loop_body_in_t_stream_t_to_slv(data : chacha20_decrypt_loop_body_in_t_stream_t) return std_logic_vector;

  function slv_to_chacha20_decrypt_loop_body_in_t_stream_t(data : std_logic_vector) return chacha20_decrypt_loop_body_in_t_stream_t;

  type uint256_t_stream_t is record
  
    data : unsigned(255 downto 0);
    valid : unsigned(0 downto 0);
  end record;
  
  constant uint256_t_stream_t_NULL : uint256_t_stream_t := (
  
    data => to_unsigned(0, 256),
    valid => to_unsigned(0, 1)
  );
  
  constant uint256_t_stream_t_SLV_LEN : integer := (
  256+1
  );
  
  function uint256_t_stream_t_to_slv(data : uint256_t_stream_t) return std_logic_vector;

  function slv_to_uint256_t_stream_t(data : std_logic_vector) return uint256_t_stream_t;

  type uint128_t_stream_t is record
  
    data : unsigned(127 downto 0);
    valid : unsigned(0 downto 0);
  end record;
  
  constant uint128_t_stream_t_NULL : uint128_t_stream_t := (
  
    data => to_unsigned(0, 128),
    valid => to_unsigned(0, 1)
  );
  
  constant uint128_t_stream_t_SLV_LEN : integer := (
  128+1
  );
  
  function uint128_t_stream_t_to_slv(data : uint128_t_stream_t) return std_logic_vector;

  function slv_to_uint128_t_stream_t(data : std_logic_vector) return uint128_t_stream_t;

  type u320_t is record
  
    limbs : uint64_t_5;
  end record;
  
  constant u320_t_NULL : u320_t := (
  
    limbs => (others => to_unsigned(0, 64))
  );
  
  constant u320_t_SLV_LEN : integer := (
  uint64_t_5_SLV_LEN
  );
  
  function u320_t_to_slv(data : u320_t) return std_logic_vector;

  function slv_to_u320_t(data : std_logic_vector) return u320_t;

  type u8_16_t is record
  
    bytes : uint8_t_16;
  end record;
  
  constant u8_16_t_NULL : u8_16_t := (
  
    bytes => (others => to_unsigned(0, 8))
  );
  
  constant u8_16_t_SLV_LEN : integer := (
  uint8_t_16_SLV_LEN
  );
  
  function u8_16_t_to_slv(data : u8_16_t) return std_logic_vector;

  function slv_to_u8_16_t(data : std_logic_vector) return u8_16_t;

  type poly1305_mac_loop_body_in_t is record
  
    block_bytes : uint8_t_16;
    r : u320_t;
    a : u320_t;
  end record;
  
  constant poly1305_mac_loop_body_in_t_NULL : poly1305_mac_loop_body_in_t := (
  
    block_bytes => (others => to_unsigned(0, 8)),
    r => u320_t_NULL,
    a => u320_t_NULL
  );
  
  constant poly1305_mac_loop_body_in_t_SLV_LEN : integer := (
  uint8_t_16_SLV_LEN+u320_t_SLV_LEN+u320_t_SLV_LEN
  );
  
  function poly1305_mac_loop_body_in_t_to_slv(data : poly1305_mac_loop_body_in_t) return std_logic_vector;

  function slv_to_poly1305_mac_loop_body_in_t(data : std_logic_vector) return poly1305_mac_loop_body_in_t;

  type chacha20_decrypt_pipeline_no_handshake_in_reg_t is record
  
    data : chacha20_decrypt_loop_body_in_t;
    id : unsigned(7 downto 0);
    valid : unsigned(0 downto 0);
  end record;
  
  constant chacha20_decrypt_pipeline_no_handshake_in_reg_t_NULL : chacha20_decrypt_pipeline_no_handshake_in_reg_t := (
  
    data => chacha20_decrypt_loop_body_in_t_NULL,
    id => to_unsigned(0, 8),
    valid => to_unsigned(0, 1)
  );
  
  constant chacha20_decrypt_pipeline_no_handshake_in_reg_t_SLV_LEN : integer := (
  chacha20_decrypt_loop_body_in_t_SLV_LEN+8+1
  );
  
  function chacha20_decrypt_pipeline_no_handshake_in_reg_t_to_slv(data : chacha20_decrypt_pipeline_no_handshake_in_reg_t) return std_logic_vector;

  function slv_to_chacha20_decrypt_pipeline_no_handshake_in_reg_t(data : std_logic_vector) return chacha20_decrypt_pipeline_no_handshake_in_reg_t;

  type chacha20_decrypt_pipeline_no_handshake_out_reg_t is record
  
    data : axis512_t;
    id : unsigned(7 downto 0);
    valid : unsigned(0 downto 0);
  end record;
  
  constant chacha20_decrypt_pipeline_no_handshake_out_reg_t_NULL : chacha20_decrypt_pipeline_no_handshake_out_reg_t := (
  
    data => axis512_t_NULL,
    id => to_unsigned(0, 8),
    valid => to_unsigned(0, 1)
  );
  
  constant chacha20_decrypt_pipeline_no_handshake_out_reg_t_SLV_LEN : integer := (
  axis512_t_SLV_LEN+8+1
  );
  
  function chacha20_decrypt_pipeline_no_handshake_out_reg_t_to_slv(data : chacha20_decrypt_pipeline_no_handshake_out_reg_t) return std_logic_vector;

  function slv_to_chacha20_decrypt_pipeline_no_handshake_out_reg_t(data : std_logic_vector) return chacha20_decrypt_pipeline_no_handshake_out_reg_t;

  type chacha20_decrypt_pipeline_FIFO_t is record
  
    data_out : axis512_t;
    data_out_valid : unsigned(0 downto 0);
    data_in_ready : unsigned(0 downto 0);
  end record;
  
  constant chacha20_decrypt_pipeline_FIFO_t_NULL : chacha20_decrypt_pipeline_FIFO_t := (
  
    data_out => axis512_t_NULL,
    data_out_valid => to_unsigned(0, 1),
    data_in_ready => to_unsigned(0, 1)
  );
  
  constant chacha20_decrypt_pipeline_FIFO_t_SLV_LEN : integer := (
  axis512_t_SLV_LEN+1+1
  );
  
  function chacha20_decrypt_pipeline_FIFO_t_to_slv(data : chacha20_decrypt_pipeline_FIFO_t) return std_logic_vector;

  function slv_to_chacha20_decrypt_pipeline_FIFO_t(data : std_logic_vector) return chacha20_decrypt_pipeline_FIFO_t;

  type poly1305_pipeline_in_reg_t is record
  
    data : poly1305_mac_loop_body_in_t;
    id : unsigned(7 downto 0);
    valid : unsigned(0 downto 0);
  end record;
  
  constant poly1305_pipeline_in_reg_t_NULL : poly1305_pipeline_in_reg_t := (
  
    data => poly1305_mac_loop_body_in_t_NULL,
    id => to_unsigned(0, 8),
    valid => to_unsigned(0, 1)
  );
  
  constant poly1305_pipeline_in_reg_t_SLV_LEN : integer := (
  poly1305_mac_loop_body_in_t_SLV_LEN+8+1
  );
  
  function poly1305_pipeline_in_reg_t_to_slv(data : poly1305_pipeline_in_reg_t) return std_logic_vector;

  function slv_to_poly1305_pipeline_in_reg_t(data : std_logic_vector) return poly1305_pipeline_in_reg_t;

  type poly1305_pipeline_out_reg_t is record
  
    data : u320_t;
    id : unsigned(7 downto 0);
    valid : unsigned(0 downto 0);
  end record;
  
  constant poly1305_pipeline_out_reg_t_NULL : poly1305_pipeline_out_reg_t := (
  
    data => u320_t_NULL,
    id => to_unsigned(0, 8),
    valid => to_unsigned(0, 1)
  );
  
  constant poly1305_pipeline_out_reg_t_SLV_LEN : integer := (
  u320_t_SLV_LEN+8+1
  );
  
  function poly1305_pipeline_out_reg_t_to_slv(data : poly1305_pipeline_out_reg_t) return std_logic_vector;

  function slv_to_poly1305_pipeline_out_reg_t(data : std_logic_vector) return poly1305_pipeline_out_reg_t;

  type uint1_t_stream_t is record
  
    data : unsigned(0 downto 0);
    valid : unsigned(0 downto 0);
  end record;
  
  constant uint1_t_stream_t_NULL : uint1_t_stream_t := (
  
    data => to_unsigned(0, 1),
    valid => to_unsigned(0, 1)
  );
  
  constant uint1_t_stream_t_SLV_LEN : integer := (
  1+1
  );
  
  function uint1_t_stream_t_to_slv(data : uint1_t_stream_t) return std_logic_vector;

  function slv_to_uint1_t_stream_t(data : std_logic_vector) return uint1_t_stream_t;

  type verify_fifo_FIFO_write_t is record
  
    ready : unsigned(0 downto 0);
  end record;
  
  constant verify_fifo_FIFO_write_t_NULL : verify_fifo_FIFO_write_t := (
  
    ready => to_unsigned(0, 1)
  );
  
  constant verify_fifo_FIFO_write_t_SLV_LEN : integer := (
  1
  );
  
  function verify_fifo_FIFO_write_t_to_slv(data : verify_fifo_FIFO_write_t) return std_logic_vector;

  function slv_to_verify_fifo_FIFO_write_t(data : std_logic_vector) return verify_fifo_FIFO_write_t;

  type uint8_t_array_64_t is record
  
    data : uint8_t_64;
  end record;
  
  constant uint8_t_array_64_t_NULL : uint8_t_array_64_t := (
  
    data => (others => to_unsigned(0, 8))
  );
  
  constant uint8_t_array_64_t_SLV_LEN : integer := (
  uint8_t_64_SLV_LEN
  );
  
  function uint8_t_array_64_t_to_slv(data : uint8_t_array_64_t) return std_logic_vector;

  function slv_to_uint8_t_array_64_t(data : std_logic_vector) return uint8_t_array_64_t;

  type uint8_t_array_40_t is record
  
    data : uint8_t_40;
  end record;
  
  constant uint8_t_array_40_t_NULL : uint8_t_array_40_t := (
  
    data => (others => to_unsigned(0, 8))
  );
  
  constant uint8_t_array_40_t_SLV_LEN : integer := (
  uint8_t_40_SLV_LEN
  );
  
  function uint8_t_array_40_t_to_slv(data : uint8_t_array_40_t) return std_logic_vector;

  function slv_to_uint8_t_array_40_t(data : std_logic_vector) return uint8_t_array_40_t;

  type uint8_t_array_8_t is record
  
    data : uint8_t_8;
  end record;
  
  constant uint8_t_array_8_t_NULL : uint8_t_array_8_t := (
  
    data => (others => to_unsigned(0, 8))
  );
  
  constant uint8_t_array_8_t_SLV_LEN : integer := (
  uint8_t_8_SLV_LEN
  );
  
  function uint8_t_array_8_t_to_slv(data : uint8_t_array_8_t) return std_logic_vector;

  function slv_to_uint8_t_array_8_t(data : std_logic_vector) return uint8_t_array_8_t;

  type uint8_t_array_4_t is record
  
    data : uint8_t_4;
  end record;
  
  constant uint8_t_array_4_t_NULL : uint8_t_array_4_t := (
  
    data => (others => to_unsigned(0, 8))
  );
  
  constant uint8_t_array_4_t_SLV_LEN : integer := (
  uint8_t_4_SLV_LEN
  );
  
  function uint8_t_array_4_t_to_slv(data : uint8_t_array_4_t) return std_logic_vector;

  function slv_to_uint8_t_array_4_t(data : std_logic_vector) return uint8_t_array_4_t;

  type uint32_t_array_16_t is record
  
    data : uint32_t_16;
  end record;
  
  constant uint32_t_array_16_t_NULL : uint32_t_array_16_t := (
  
    data => (others => to_unsigned(0, 32))
  );
  
  constant uint32_t_array_16_t_SLV_LEN : integer := (
  uint32_t_16_SLV_LEN
  );
  
  function uint32_t_array_16_t_to_slv(data : uint32_t_array_16_t) return std_logic_vector;

  function slv_to_uint32_t_array_16_t(data : std_logic_vector) return uint32_t_array_16_t;

  type uint8_t_array_144_t is record
  
    data : uint8_t_144;
  end record;
  
  constant uint8_t_array_144_t_NULL : uint8_t_array_144_t := (
  
    data => (others => to_unsigned(0, 8))
  );
  
  constant uint8_t_array_144_t_SLV_LEN : integer := (
  uint8_t_144_SLV_LEN
  );
  
  function uint8_t_array_144_t_to_slv(data : uint8_t_array_144_t) return std_logic_vector;

  function slv_to_uint8_t_array_144_t(data : std_logic_vector) return uint8_t_array_144_t;

  type char_array_128_t is record
  
    data : char_128;
  end record;
  
  constant char_array_128_t_NULL : char_array_128_t := (
  
    data => (others => to_unsigned(0, 8))
  );
  
  constant char_array_128_t_SLV_LEN : integer := (
  char_128_SLV_LEN
  );
  
  function char_array_128_t_to_slv(data : char_array_128_t) return std_logic_vector;

  function slv_to_char_array_128_t(data : std_logic_vector) return char_array_128_t;
type axis128_t_stream_t_4 is array(0 to 3) of axis128_t_stream_t;
constant axis128_t_stream_t_4_SLV_LEN : integer := axis128_t_stream_t_SLV_LEN * 4;

      function axis128_t_stream_t_4_to_slv(data : axis128_t_stream_t_4) return std_logic_vector;

      function slv_to_axis128_t_stream_t_4(data : std_logic_vector) return axis128_t_stream_t_4;
type axis128_t_1 is array(0 to 0) of axis128_t;
constant axis128_t_1_SLV_LEN : integer := axis128_t_SLV_LEN * 1;

      function axis128_t_1_to_slv(data : axis128_t_1) return std_logic_vector;

      function slv_to_axis128_t_1(data : std_logic_vector) return axis128_t_1;

  type axis512_to_axis128_array_t is record
  
    axis_chunks : axis128_t_stream_t_4;
  end record;
  
  constant axis512_to_axis128_array_t_NULL : axis512_to_axis128_array_t := (
  
    axis_chunks => (others => axis128_t_stream_t_NULL)
  );
  
  constant axis512_to_axis128_array_t_SLV_LEN : integer := (
  axis128_t_stream_t_4_SLV_LEN
  );
  
  function axis512_to_axis128_array_t_to_slv(data : axis512_to_axis128_array_t) return std_logic_vector;

  function slv_to_axis512_to_axis128_array_t(data : std_logic_vector) return axis512_to_axis128_array_t;

  type verify_fifo_FIFO_read_t is record
  
    data : axis128_t_1;
    valid : unsigned(0 downto 0);
  end record;
  
  constant verify_fifo_FIFO_read_t_NULL : verify_fifo_FIFO_read_t := (
  
    data => (others => axis128_t_NULL),
    valid => to_unsigned(0, 1)
  );
  
  constant verify_fifo_FIFO_read_t_SLV_LEN : integer := (
  axis128_t_1_SLV_LEN+1
  );
  
  function verify_fifo_FIFO_read_t_to_slv(data : verify_fifo_FIFO_read_t) return std_logic_vector;

  function slv_to_verify_fifo_FIFO_read_t(data : std_logic_vector) return verify_fifo_FIFO_read_t;

end c_structs_pkg;
package body c_structs_pkg is
function uint1_t_to_slv(x : uint1_t) return std_logic_vector is
  variable rv : std_logic_vector(0 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1_t(x : std_logic_vector) return uint1_t is
  variable rv : uint1_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function uint2_t_to_slv(x : uint2_t) return std_logic_vector is
  variable rv : std_logic_vector(1 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2_t(x : std_logic_vector) return uint2_t is
  variable rv : uint2_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2_t_to_slv(x : int2_t) return std_logic_vector is
  variable rv : std_logic_vector(1 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2_t(x : std_logic_vector) return int2_t is
  variable rv : int2_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint3_t_to_slv(x : uint3_t) return std_logic_vector is
  variable rv : std_logic_vector(2 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint3_t(x : std_logic_vector) return uint3_t is
  variable rv : uint3_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int3_t_to_slv(x : int3_t) return std_logic_vector is
  variable rv : std_logic_vector(2 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int3_t(x : std_logic_vector) return int3_t is
  variable rv : int3_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint4_t_to_slv(x : uint4_t) return std_logic_vector is
  variable rv : std_logic_vector(3 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint4_t(x : std_logic_vector) return uint4_t is
  variable rv : uint4_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int4_t_to_slv(x : int4_t) return std_logic_vector is
  variable rv : std_logic_vector(3 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int4_t(x : std_logic_vector) return int4_t is
  variable rv : int4_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint5_t_to_slv(x : uint5_t) return std_logic_vector is
  variable rv : std_logic_vector(4 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint5_t(x : std_logic_vector) return uint5_t is
  variable rv : uint5_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int5_t_to_slv(x : int5_t) return std_logic_vector is
  variable rv : std_logic_vector(4 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int5_t(x : std_logic_vector) return int5_t is
  variable rv : int5_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint6_t_to_slv(x : uint6_t) return std_logic_vector is
  variable rv : std_logic_vector(5 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint6_t(x : std_logic_vector) return uint6_t is
  variable rv : uint6_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int6_t_to_slv(x : int6_t) return std_logic_vector is
  variable rv : std_logic_vector(5 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int6_t(x : std_logic_vector) return int6_t is
  variable rv : int6_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint7_t_to_slv(x : uint7_t) return std_logic_vector is
  variable rv : std_logic_vector(6 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint7_t(x : std_logic_vector) return uint7_t is
  variable rv : uint7_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int7_t_to_slv(x : int7_t) return std_logic_vector is
  variable rv : std_logic_vector(6 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int7_t(x : std_logic_vector) return int7_t is
  variable rv : int7_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint8_t_to_slv(x : uint8_t) return std_logic_vector is
  variable rv : std_logic_vector(7 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint8_t(x : std_logic_vector) return uint8_t is
  variable rv : uint8_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int8_t_to_slv(x : int8_t) return std_logic_vector is
  variable rv : std_logic_vector(7 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int8_t(x : std_logic_vector) return int8_t is
  variable rv : int8_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint9_t_to_slv(x : uint9_t) return std_logic_vector is
  variable rv : std_logic_vector(8 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint9_t(x : std_logic_vector) return uint9_t is
  variable rv : uint9_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int9_t_to_slv(x : int9_t) return std_logic_vector is
  variable rv : std_logic_vector(8 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int9_t(x : std_logic_vector) return int9_t is
  variable rv : int9_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint10_t_to_slv(x : uint10_t) return std_logic_vector is
  variable rv : std_logic_vector(9 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint10_t(x : std_logic_vector) return uint10_t is
  variable rv : uint10_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int10_t_to_slv(x : int10_t) return std_logic_vector is
  variable rv : std_logic_vector(9 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int10_t(x : std_logic_vector) return int10_t is
  variable rv : int10_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint11_t_to_slv(x : uint11_t) return std_logic_vector is
  variable rv : std_logic_vector(10 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint11_t(x : std_logic_vector) return uint11_t is
  variable rv : uint11_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int11_t_to_slv(x : int11_t) return std_logic_vector is
  variable rv : std_logic_vector(10 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int11_t(x : std_logic_vector) return int11_t is
  variable rv : int11_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint12_t_to_slv(x : uint12_t) return std_logic_vector is
  variable rv : std_logic_vector(11 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint12_t(x : std_logic_vector) return uint12_t is
  variable rv : uint12_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int12_t_to_slv(x : int12_t) return std_logic_vector is
  variable rv : std_logic_vector(11 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int12_t(x : std_logic_vector) return int12_t is
  variable rv : int12_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint13_t_to_slv(x : uint13_t) return std_logic_vector is
  variable rv : std_logic_vector(12 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint13_t(x : std_logic_vector) return uint13_t is
  variable rv : uint13_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int13_t_to_slv(x : int13_t) return std_logic_vector is
  variable rv : std_logic_vector(12 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int13_t(x : std_logic_vector) return int13_t is
  variable rv : int13_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint14_t_to_slv(x : uint14_t) return std_logic_vector is
  variable rv : std_logic_vector(13 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint14_t(x : std_logic_vector) return uint14_t is
  variable rv : uint14_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int14_t_to_slv(x : int14_t) return std_logic_vector is
  variable rv : std_logic_vector(13 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int14_t(x : std_logic_vector) return int14_t is
  variable rv : int14_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint15_t_to_slv(x : uint15_t) return std_logic_vector is
  variable rv : std_logic_vector(14 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint15_t(x : std_logic_vector) return uint15_t is
  variable rv : uint15_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int15_t_to_slv(x : int15_t) return std_logic_vector is
  variable rv : std_logic_vector(14 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int15_t(x : std_logic_vector) return int15_t is
  variable rv : int15_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint16_t_to_slv(x : uint16_t) return std_logic_vector is
  variable rv : std_logic_vector(15 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint16_t(x : std_logic_vector) return uint16_t is
  variable rv : uint16_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int16_t_to_slv(x : int16_t) return std_logic_vector is
  variable rv : std_logic_vector(15 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int16_t(x : std_logic_vector) return int16_t is
  variable rv : int16_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint17_t_to_slv(x : uint17_t) return std_logic_vector is
  variable rv : std_logic_vector(16 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint17_t(x : std_logic_vector) return uint17_t is
  variable rv : uint17_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int17_t_to_slv(x : int17_t) return std_logic_vector is
  variable rv : std_logic_vector(16 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int17_t(x : std_logic_vector) return int17_t is
  variable rv : int17_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint18_t_to_slv(x : uint18_t) return std_logic_vector is
  variable rv : std_logic_vector(17 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint18_t(x : std_logic_vector) return uint18_t is
  variable rv : uint18_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int18_t_to_slv(x : int18_t) return std_logic_vector is
  variable rv : std_logic_vector(17 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int18_t(x : std_logic_vector) return int18_t is
  variable rv : int18_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint19_t_to_slv(x : uint19_t) return std_logic_vector is
  variable rv : std_logic_vector(18 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint19_t(x : std_logic_vector) return uint19_t is
  variable rv : uint19_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int19_t_to_slv(x : int19_t) return std_logic_vector is
  variable rv : std_logic_vector(18 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int19_t(x : std_logic_vector) return int19_t is
  variable rv : int19_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint20_t_to_slv(x : uint20_t) return std_logic_vector is
  variable rv : std_logic_vector(19 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint20_t(x : std_logic_vector) return uint20_t is
  variable rv : uint20_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int20_t_to_slv(x : int20_t) return std_logic_vector is
  variable rv : std_logic_vector(19 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int20_t(x : std_logic_vector) return int20_t is
  variable rv : int20_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint21_t_to_slv(x : uint21_t) return std_logic_vector is
  variable rv : std_logic_vector(20 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint21_t(x : std_logic_vector) return uint21_t is
  variable rv : uint21_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int21_t_to_slv(x : int21_t) return std_logic_vector is
  variable rv : std_logic_vector(20 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int21_t(x : std_logic_vector) return int21_t is
  variable rv : int21_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint22_t_to_slv(x : uint22_t) return std_logic_vector is
  variable rv : std_logic_vector(21 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint22_t(x : std_logic_vector) return uint22_t is
  variable rv : uint22_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int22_t_to_slv(x : int22_t) return std_logic_vector is
  variable rv : std_logic_vector(21 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int22_t(x : std_logic_vector) return int22_t is
  variable rv : int22_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint23_t_to_slv(x : uint23_t) return std_logic_vector is
  variable rv : std_logic_vector(22 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint23_t(x : std_logic_vector) return uint23_t is
  variable rv : uint23_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int23_t_to_slv(x : int23_t) return std_logic_vector is
  variable rv : std_logic_vector(22 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int23_t(x : std_logic_vector) return int23_t is
  variable rv : int23_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint24_t_to_slv(x : uint24_t) return std_logic_vector is
  variable rv : std_logic_vector(23 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint24_t(x : std_logic_vector) return uint24_t is
  variable rv : uint24_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int24_t_to_slv(x : int24_t) return std_logic_vector is
  variable rv : std_logic_vector(23 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int24_t(x : std_logic_vector) return int24_t is
  variable rv : int24_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint25_t_to_slv(x : uint25_t) return std_logic_vector is
  variable rv : std_logic_vector(24 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint25_t(x : std_logic_vector) return uint25_t is
  variable rv : uint25_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int25_t_to_slv(x : int25_t) return std_logic_vector is
  variable rv : std_logic_vector(24 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int25_t(x : std_logic_vector) return int25_t is
  variable rv : int25_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint26_t_to_slv(x : uint26_t) return std_logic_vector is
  variable rv : std_logic_vector(25 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint26_t(x : std_logic_vector) return uint26_t is
  variable rv : uint26_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int26_t_to_slv(x : int26_t) return std_logic_vector is
  variable rv : std_logic_vector(25 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int26_t(x : std_logic_vector) return int26_t is
  variable rv : int26_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint27_t_to_slv(x : uint27_t) return std_logic_vector is
  variable rv : std_logic_vector(26 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint27_t(x : std_logic_vector) return uint27_t is
  variable rv : uint27_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int27_t_to_slv(x : int27_t) return std_logic_vector is
  variable rv : std_logic_vector(26 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int27_t(x : std_logic_vector) return int27_t is
  variable rv : int27_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint28_t_to_slv(x : uint28_t) return std_logic_vector is
  variable rv : std_logic_vector(27 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint28_t(x : std_logic_vector) return uint28_t is
  variable rv : uint28_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int28_t_to_slv(x : int28_t) return std_logic_vector is
  variable rv : std_logic_vector(27 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int28_t(x : std_logic_vector) return int28_t is
  variable rv : int28_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint29_t_to_slv(x : uint29_t) return std_logic_vector is
  variable rv : std_logic_vector(28 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint29_t(x : std_logic_vector) return uint29_t is
  variable rv : uint29_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int29_t_to_slv(x : int29_t) return std_logic_vector is
  variable rv : std_logic_vector(28 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int29_t(x : std_logic_vector) return int29_t is
  variable rv : int29_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint30_t_to_slv(x : uint30_t) return std_logic_vector is
  variable rv : std_logic_vector(29 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint30_t(x : std_logic_vector) return uint30_t is
  variable rv : uint30_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int30_t_to_slv(x : int30_t) return std_logic_vector is
  variable rv : std_logic_vector(29 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int30_t(x : std_logic_vector) return int30_t is
  variable rv : int30_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint31_t_to_slv(x : uint31_t) return std_logic_vector is
  variable rv : std_logic_vector(30 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint31_t(x : std_logic_vector) return uint31_t is
  variable rv : uint31_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int31_t_to_slv(x : int31_t) return std_logic_vector is
  variable rv : std_logic_vector(30 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int31_t(x : std_logic_vector) return int31_t is
  variable rv : int31_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint32_t_to_slv(x : uint32_t) return std_logic_vector is
  variable rv : std_logic_vector(31 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint32_t(x : std_logic_vector) return uint32_t is
  variable rv : uint32_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int32_t_to_slv(x : int32_t) return std_logic_vector is
  variable rv : std_logic_vector(31 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int32_t(x : std_logic_vector) return int32_t is
  variable rv : int32_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint33_t_to_slv(x : uint33_t) return std_logic_vector is
  variable rv : std_logic_vector(32 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint33_t(x : std_logic_vector) return uint33_t is
  variable rv : uint33_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int33_t_to_slv(x : int33_t) return std_logic_vector is
  variable rv : std_logic_vector(32 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int33_t(x : std_logic_vector) return int33_t is
  variable rv : int33_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint34_t_to_slv(x : uint34_t) return std_logic_vector is
  variable rv : std_logic_vector(33 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint34_t(x : std_logic_vector) return uint34_t is
  variable rv : uint34_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int34_t_to_slv(x : int34_t) return std_logic_vector is
  variable rv : std_logic_vector(33 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int34_t(x : std_logic_vector) return int34_t is
  variable rv : int34_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint35_t_to_slv(x : uint35_t) return std_logic_vector is
  variable rv : std_logic_vector(34 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint35_t(x : std_logic_vector) return uint35_t is
  variable rv : uint35_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int35_t_to_slv(x : int35_t) return std_logic_vector is
  variable rv : std_logic_vector(34 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int35_t(x : std_logic_vector) return int35_t is
  variable rv : int35_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint36_t_to_slv(x : uint36_t) return std_logic_vector is
  variable rv : std_logic_vector(35 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint36_t(x : std_logic_vector) return uint36_t is
  variable rv : uint36_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int36_t_to_slv(x : int36_t) return std_logic_vector is
  variable rv : std_logic_vector(35 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int36_t(x : std_logic_vector) return int36_t is
  variable rv : int36_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint37_t_to_slv(x : uint37_t) return std_logic_vector is
  variable rv : std_logic_vector(36 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint37_t(x : std_logic_vector) return uint37_t is
  variable rv : uint37_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int37_t_to_slv(x : int37_t) return std_logic_vector is
  variable rv : std_logic_vector(36 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int37_t(x : std_logic_vector) return int37_t is
  variable rv : int37_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint38_t_to_slv(x : uint38_t) return std_logic_vector is
  variable rv : std_logic_vector(37 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint38_t(x : std_logic_vector) return uint38_t is
  variable rv : uint38_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int38_t_to_slv(x : int38_t) return std_logic_vector is
  variable rv : std_logic_vector(37 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int38_t(x : std_logic_vector) return int38_t is
  variable rv : int38_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint39_t_to_slv(x : uint39_t) return std_logic_vector is
  variable rv : std_logic_vector(38 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint39_t(x : std_logic_vector) return uint39_t is
  variable rv : uint39_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int39_t_to_slv(x : int39_t) return std_logic_vector is
  variable rv : std_logic_vector(38 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int39_t(x : std_logic_vector) return int39_t is
  variable rv : int39_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint40_t_to_slv(x : uint40_t) return std_logic_vector is
  variable rv : std_logic_vector(39 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint40_t(x : std_logic_vector) return uint40_t is
  variable rv : uint40_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int40_t_to_slv(x : int40_t) return std_logic_vector is
  variable rv : std_logic_vector(39 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int40_t(x : std_logic_vector) return int40_t is
  variable rv : int40_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint41_t_to_slv(x : uint41_t) return std_logic_vector is
  variable rv : std_logic_vector(40 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint41_t(x : std_logic_vector) return uint41_t is
  variable rv : uint41_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int41_t_to_slv(x : int41_t) return std_logic_vector is
  variable rv : std_logic_vector(40 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int41_t(x : std_logic_vector) return int41_t is
  variable rv : int41_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint42_t_to_slv(x : uint42_t) return std_logic_vector is
  variable rv : std_logic_vector(41 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint42_t(x : std_logic_vector) return uint42_t is
  variable rv : uint42_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int42_t_to_slv(x : int42_t) return std_logic_vector is
  variable rv : std_logic_vector(41 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int42_t(x : std_logic_vector) return int42_t is
  variable rv : int42_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint43_t_to_slv(x : uint43_t) return std_logic_vector is
  variable rv : std_logic_vector(42 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint43_t(x : std_logic_vector) return uint43_t is
  variable rv : uint43_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int43_t_to_slv(x : int43_t) return std_logic_vector is
  variable rv : std_logic_vector(42 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int43_t(x : std_logic_vector) return int43_t is
  variable rv : int43_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint44_t_to_slv(x : uint44_t) return std_logic_vector is
  variable rv : std_logic_vector(43 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint44_t(x : std_logic_vector) return uint44_t is
  variable rv : uint44_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int44_t_to_slv(x : int44_t) return std_logic_vector is
  variable rv : std_logic_vector(43 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int44_t(x : std_logic_vector) return int44_t is
  variable rv : int44_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint45_t_to_slv(x : uint45_t) return std_logic_vector is
  variable rv : std_logic_vector(44 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint45_t(x : std_logic_vector) return uint45_t is
  variable rv : uint45_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int45_t_to_slv(x : int45_t) return std_logic_vector is
  variable rv : std_logic_vector(44 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int45_t(x : std_logic_vector) return int45_t is
  variable rv : int45_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint46_t_to_slv(x : uint46_t) return std_logic_vector is
  variable rv : std_logic_vector(45 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint46_t(x : std_logic_vector) return uint46_t is
  variable rv : uint46_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int46_t_to_slv(x : int46_t) return std_logic_vector is
  variable rv : std_logic_vector(45 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int46_t(x : std_logic_vector) return int46_t is
  variable rv : int46_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint47_t_to_slv(x : uint47_t) return std_logic_vector is
  variable rv : std_logic_vector(46 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint47_t(x : std_logic_vector) return uint47_t is
  variable rv : uint47_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int47_t_to_slv(x : int47_t) return std_logic_vector is
  variable rv : std_logic_vector(46 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int47_t(x : std_logic_vector) return int47_t is
  variable rv : int47_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint48_t_to_slv(x : uint48_t) return std_logic_vector is
  variable rv : std_logic_vector(47 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint48_t(x : std_logic_vector) return uint48_t is
  variable rv : uint48_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int48_t_to_slv(x : int48_t) return std_logic_vector is
  variable rv : std_logic_vector(47 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int48_t(x : std_logic_vector) return int48_t is
  variable rv : int48_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint49_t_to_slv(x : uint49_t) return std_logic_vector is
  variable rv : std_logic_vector(48 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint49_t(x : std_logic_vector) return uint49_t is
  variable rv : uint49_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int49_t_to_slv(x : int49_t) return std_logic_vector is
  variable rv : std_logic_vector(48 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int49_t(x : std_logic_vector) return int49_t is
  variable rv : int49_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint50_t_to_slv(x : uint50_t) return std_logic_vector is
  variable rv : std_logic_vector(49 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint50_t(x : std_logic_vector) return uint50_t is
  variable rv : uint50_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int50_t_to_slv(x : int50_t) return std_logic_vector is
  variable rv : std_logic_vector(49 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int50_t(x : std_logic_vector) return int50_t is
  variable rv : int50_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint51_t_to_slv(x : uint51_t) return std_logic_vector is
  variable rv : std_logic_vector(50 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint51_t(x : std_logic_vector) return uint51_t is
  variable rv : uint51_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int51_t_to_slv(x : int51_t) return std_logic_vector is
  variable rv : std_logic_vector(50 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int51_t(x : std_logic_vector) return int51_t is
  variable rv : int51_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint52_t_to_slv(x : uint52_t) return std_logic_vector is
  variable rv : std_logic_vector(51 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint52_t(x : std_logic_vector) return uint52_t is
  variable rv : uint52_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int52_t_to_slv(x : int52_t) return std_logic_vector is
  variable rv : std_logic_vector(51 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int52_t(x : std_logic_vector) return int52_t is
  variable rv : int52_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint53_t_to_slv(x : uint53_t) return std_logic_vector is
  variable rv : std_logic_vector(52 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint53_t(x : std_logic_vector) return uint53_t is
  variable rv : uint53_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int53_t_to_slv(x : int53_t) return std_logic_vector is
  variable rv : std_logic_vector(52 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int53_t(x : std_logic_vector) return int53_t is
  variable rv : int53_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint54_t_to_slv(x : uint54_t) return std_logic_vector is
  variable rv : std_logic_vector(53 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint54_t(x : std_logic_vector) return uint54_t is
  variable rv : uint54_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int54_t_to_slv(x : int54_t) return std_logic_vector is
  variable rv : std_logic_vector(53 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int54_t(x : std_logic_vector) return int54_t is
  variable rv : int54_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint55_t_to_slv(x : uint55_t) return std_logic_vector is
  variable rv : std_logic_vector(54 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint55_t(x : std_logic_vector) return uint55_t is
  variable rv : uint55_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int55_t_to_slv(x : int55_t) return std_logic_vector is
  variable rv : std_logic_vector(54 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int55_t(x : std_logic_vector) return int55_t is
  variable rv : int55_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint56_t_to_slv(x : uint56_t) return std_logic_vector is
  variable rv : std_logic_vector(55 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint56_t(x : std_logic_vector) return uint56_t is
  variable rv : uint56_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int56_t_to_slv(x : int56_t) return std_logic_vector is
  variable rv : std_logic_vector(55 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int56_t(x : std_logic_vector) return int56_t is
  variable rv : int56_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint57_t_to_slv(x : uint57_t) return std_logic_vector is
  variable rv : std_logic_vector(56 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint57_t(x : std_logic_vector) return uint57_t is
  variable rv : uint57_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int57_t_to_slv(x : int57_t) return std_logic_vector is
  variable rv : std_logic_vector(56 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int57_t(x : std_logic_vector) return int57_t is
  variable rv : int57_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint58_t_to_slv(x : uint58_t) return std_logic_vector is
  variable rv : std_logic_vector(57 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint58_t(x : std_logic_vector) return uint58_t is
  variable rv : uint58_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int58_t_to_slv(x : int58_t) return std_logic_vector is
  variable rv : std_logic_vector(57 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int58_t(x : std_logic_vector) return int58_t is
  variable rv : int58_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint59_t_to_slv(x : uint59_t) return std_logic_vector is
  variable rv : std_logic_vector(58 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint59_t(x : std_logic_vector) return uint59_t is
  variable rv : uint59_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int59_t_to_slv(x : int59_t) return std_logic_vector is
  variable rv : std_logic_vector(58 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int59_t(x : std_logic_vector) return int59_t is
  variable rv : int59_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint60_t_to_slv(x : uint60_t) return std_logic_vector is
  variable rv : std_logic_vector(59 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint60_t(x : std_logic_vector) return uint60_t is
  variable rv : uint60_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int60_t_to_slv(x : int60_t) return std_logic_vector is
  variable rv : std_logic_vector(59 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int60_t(x : std_logic_vector) return int60_t is
  variable rv : int60_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint61_t_to_slv(x : uint61_t) return std_logic_vector is
  variable rv : std_logic_vector(60 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint61_t(x : std_logic_vector) return uint61_t is
  variable rv : uint61_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int61_t_to_slv(x : int61_t) return std_logic_vector is
  variable rv : std_logic_vector(60 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int61_t(x : std_logic_vector) return int61_t is
  variable rv : int61_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint62_t_to_slv(x : uint62_t) return std_logic_vector is
  variable rv : std_logic_vector(61 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint62_t(x : std_logic_vector) return uint62_t is
  variable rv : uint62_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int62_t_to_slv(x : int62_t) return std_logic_vector is
  variable rv : std_logic_vector(61 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int62_t(x : std_logic_vector) return int62_t is
  variable rv : int62_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint63_t_to_slv(x : uint63_t) return std_logic_vector is
  variable rv : std_logic_vector(62 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint63_t(x : std_logic_vector) return uint63_t is
  variable rv : uint63_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int63_t_to_slv(x : int63_t) return std_logic_vector is
  variable rv : std_logic_vector(62 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int63_t(x : std_logic_vector) return int63_t is
  variable rv : int63_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint64_t_to_slv(x : uint64_t) return std_logic_vector is
  variable rv : std_logic_vector(63 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint64_t(x : std_logic_vector) return uint64_t is
  variable rv : uint64_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int64_t_to_slv(x : int64_t) return std_logic_vector is
  variable rv : std_logic_vector(63 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int64_t(x : std_logic_vector) return int64_t is
  variable rv : int64_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint65_t_to_slv(x : uint65_t) return std_logic_vector is
  variable rv : std_logic_vector(64 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint65_t(x : std_logic_vector) return uint65_t is
  variable rv : uint65_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int65_t_to_slv(x : int65_t) return std_logic_vector is
  variable rv : std_logic_vector(64 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int65_t(x : std_logic_vector) return int65_t is
  variable rv : int65_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint66_t_to_slv(x : uint66_t) return std_logic_vector is
  variable rv : std_logic_vector(65 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint66_t(x : std_logic_vector) return uint66_t is
  variable rv : uint66_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int66_t_to_slv(x : int66_t) return std_logic_vector is
  variable rv : std_logic_vector(65 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int66_t(x : std_logic_vector) return int66_t is
  variable rv : int66_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint67_t_to_slv(x : uint67_t) return std_logic_vector is
  variable rv : std_logic_vector(66 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint67_t(x : std_logic_vector) return uint67_t is
  variable rv : uint67_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int67_t_to_slv(x : int67_t) return std_logic_vector is
  variable rv : std_logic_vector(66 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int67_t(x : std_logic_vector) return int67_t is
  variable rv : int67_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint68_t_to_slv(x : uint68_t) return std_logic_vector is
  variable rv : std_logic_vector(67 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint68_t(x : std_logic_vector) return uint68_t is
  variable rv : uint68_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int68_t_to_slv(x : int68_t) return std_logic_vector is
  variable rv : std_logic_vector(67 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int68_t(x : std_logic_vector) return int68_t is
  variable rv : int68_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint69_t_to_slv(x : uint69_t) return std_logic_vector is
  variable rv : std_logic_vector(68 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint69_t(x : std_logic_vector) return uint69_t is
  variable rv : uint69_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int69_t_to_slv(x : int69_t) return std_logic_vector is
  variable rv : std_logic_vector(68 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int69_t(x : std_logic_vector) return int69_t is
  variable rv : int69_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint70_t_to_slv(x : uint70_t) return std_logic_vector is
  variable rv : std_logic_vector(69 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint70_t(x : std_logic_vector) return uint70_t is
  variable rv : uint70_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int70_t_to_slv(x : int70_t) return std_logic_vector is
  variable rv : std_logic_vector(69 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int70_t(x : std_logic_vector) return int70_t is
  variable rv : int70_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint71_t_to_slv(x : uint71_t) return std_logic_vector is
  variable rv : std_logic_vector(70 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint71_t(x : std_logic_vector) return uint71_t is
  variable rv : uint71_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int71_t_to_slv(x : int71_t) return std_logic_vector is
  variable rv : std_logic_vector(70 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int71_t(x : std_logic_vector) return int71_t is
  variable rv : int71_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint72_t_to_slv(x : uint72_t) return std_logic_vector is
  variable rv : std_logic_vector(71 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint72_t(x : std_logic_vector) return uint72_t is
  variable rv : uint72_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int72_t_to_slv(x : int72_t) return std_logic_vector is
  variable rv : std_logic_vector(71 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int72_t(x : std_logic_vector) return int72_t is
  variable rv : int72_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint73_t_to_slv(x : uint73_t) return std_logic_vector is
  variable rv : std_logic_vector(72 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint73_t(x : std_logic_vector) return uint73_t is
  variable rv : uint73_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int73_t_to_slv(x : int73_t) return std_logic_vector is
  variable rv : std_logic_vector(72 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int73_t(x : std_logic_vector) return int73_t is
  variable rv : int73_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint74_t_to_slv(x : uint74_t) return std_logic_vector is
  variable rv : std_logic_vector(73 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint74_t(x : std_logic_vector) return uint74_t is
  variable rv : uint74_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int74_t_to_slv(x : int74_t) return std_logic_vector is
  variable rv : std_logic_vector(73 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int74_t(x : std_logic_vector) return int74_t is
  variable rv : int74_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint75_t_to_slv(x : uint75_t) return std_logic_vector is
  variable rv : std_logic_vector(74 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint75_t(x : std_logic_vector) return uint75_t is
  variable rv : uint75_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int75_t_to_slv(x : int75_t) return std_logic_vector is
  variable rv : std_logic_vector(74 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int75_t(x : std_logic_vector) return int75_t is
  variable rv : int75_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint76_t_to_slv(x : uint76_t) return std_logic_vector is
  variable rv : std_logic_vector(75 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint76_t(x : std_logic_vector) return uint76_t is
  variable rv : uint76_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int76_t_to_slv(x : int76_t) return std_logic_vector is
  variable rv : std_logic_vector(75 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int76_t(x : std_logic_vector) return int76_t is
  variable rv : int76_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint77_t_to_slv(x : uint77_t) return std_logic_vector is
  variable rv : std_logic_vector(76 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint77_t(x : std_logic_vector) return uint77_t is
  variable rv : uint77_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int77_t_to_slv(x : int77_t) return std_logic_vector is
  variable rv : std_logic_vector(76 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int77_t(x : std_logic_vector) return int77_t is
  variable rv : int77_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint78_t_to_slv(x : uint78_t) return std_logic_vector is
  variable rv : std_logic_vector(77 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint78_t(x : std_logic_vector) return uint78_t is
  variable rv : uint78_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int78_t_to_slv(x : int78_t) return std_logic_vector is
  variable rv : std_logic_vector(77 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int78_t(x : std_logic_vector) return int78_t is
  variable rv : int78_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint79_t_to_slv(x : uint79_t) return std_logic_vector is
  variable rv : std_logic_vector(78 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint79_t(x : std_logic_vector) return uint79_t is
  variable rv : uint79_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int79_t_to_slv(x : int79_t) return std_logic_vector is
  variable rv : std_logic_vector(78 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int79_t(x : std_logic_vector) return int79_t is
  variable rv : int79_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint80_t_to_slv(x : uint80_t) return std_logic_vector is
  variable rv : std_logic_vector(79 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint80_t(x : std_logic_vector) return uint80_t is
  variable rv : uint80_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int80_t_to_slv(x : int80_t) return std_logic_vector is
  variable rv : std_logic_vector(79 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int80_t(x : std_logic_vector) return int80_t is
  variable rv : int80_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint81_t_to_slv(x : uint81_t) return std_logic_vector is
  variable rv : std_logic_vector(80 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint81_t(x : std_logic_vector) return uint81_t is
  variable rv : uint81_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int81_t_to_slv(x : int81_t) return std_logic_vector is
  variable rv : std_logic_vector(80 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int81_t(x : std_logic_vector) return int81_t is
  variable rv : int81_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint82_t_to_slv(x : uint82_t) return std_logic_vector is
  variable rv : std_logic_vector(81 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint82_t(x : std_logic_vector) return uint82_t is
  variable rv : uint82_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int82_t_to_slv(x : int82_t) return std_logic_vector is
  variable rv : std_logic_vector(81 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int82_t(x : std_logic_vector) return int82_t is
  variable rv : int82_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint83_t_to_slv(x : uint83_t) return std_logic_vector is
  variable rv : std_logic_vector(82 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint83_t(x : std_logic_vector) return uint83_t is
  variable rv : uint83_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int83_t_to_slv(x : int83_t) return std_logic_vector is
  variable rv : std_logic_vector(82 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int83_t(x : std_logic_vector) return int83_t is
  variable rv : int83_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint84_t_to_slv(x : uint84_t) return std_logic_vector is
  variable rv : std_logic_vector(83 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint84_t(x : std_logic_vector) return uint84_t is
  variable rv : uint84_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int84_t_to_slv(x : int84_t) return std_logic_vector is
  variable rv : std_logic_vector(83 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int84_t(x : std_logic_vector) return int84_t is
  variable rv : int84_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint85_t_to_slv(x : uint85_t) return std_logic_vector is
  variable rv : std_logic_vector(84 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint85_t(x : std_logic_vector) return uint85_t is
  variable rv : uint85_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int85_t_to_slv(x : int85_t) return std_logic_vector is
  variable rv : std_logic_vector(84 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int85_t(x : std_logic_vector) return int85_t is
  variable rv : int85_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint86_t_to_slv(x : uint86_t) return std_logic_vector is
  variable rv : std_logic_vector(85 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint86_t(x : std_logic_vector) return uint86_t is
  variable rv : uint86_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int86_t_to_slv(x : int86_t) return std_logic_vector is
  variable rv : std_logic_vector(85 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int86_t(x : std_logic_vector) return int86_t is
  variable rv : int86_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint87_t_to_slv(x : uint87_t) return std_logic_vector is
  variable rv : std_logic_vector(86 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint87_t(x : std_logic_vector) return uint87_t is
  variable rv : uint87_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int87_t_to_slv(x : int87_t) return std_logic_vector is
  variable rv : std_logic_vector(86 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int87_t(x : std_logic_vector) return int87_t is
  variable rv : int87_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint88_t_to_slv(x : uint88_t) return std_logic_vector is
  variable rv : std_logic_vector(87 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint88_t(x : std_logic_vector) return uint88_t is
  variable rv : uint88_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int88_t_to_slv(x : int88_t) return std_logic_vector is
  variable rv : std_logic_vector(87 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int88_t(x : std_logic_vector) return int88_t is
  variable rv : int88_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint89_t_to_slv(x : uint89_t) return std_logic_vector is
  variable rv : std_logic_vector(88 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint89_t(x : std_logic_vector) return uint89_t is
  variable rv : uint89_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int89_t_to_slv(x : int89_t) return std_logic_vector is
  variable rv : std_logic_vector(88 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int89_t(x : std_logic_vector) return int89_t is
  variable rv : int89_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint90_t_to_slv(x : uint90_t) return std_logic_vector is
  variable rv : std_logic_vector(89 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint90_t(x : std_logic_vector) return uint90_t is
  variable rv : uint90_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int90_t_to_slv(x : int90_t) return std_logic_vector is
  variable rv : std_logic_vector(89 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int90_t(x : std_logic_vector) return int90_t is
  variable rv : int90_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint91_t_to_slv(x : uint91_t) return std_logic_vector is
  variable rv : std_logic_vector(90 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint91_t(x : std_logic_vector) return uint91_t is
  variable rv : uint91_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int91_t_to_slv(x : int91_t) return std_logic_vector is
  variable rv : std_logic_vector(90 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int91_t(x : std_logic_vector) return int91_t is
  variable rv : int91_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint92_t_to_slv(x : uint92_t) return std_logic_vector is
  variable rv : std_logic_vector(91 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint92_t(x : std_logic_vector) return uint92_t is
  variable rv : uint92_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int92_t_to_slv(x : int92_t) return std_logic_vector is
  variable rv : std_logic_vector(91 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int92_t(x : std_logic_vector) return int92_t is
  variable rv : int92_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint93_t_to_slv(x : uint93_t) return std_logic_vector is
  variable rv : std_logic_vector(92 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint93_t(x : std_logic_vector) return uint93_t is
  variable rv : uint93_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int93_t_to_slv(x : int93_t) return std_logic_vector is
  variable rv : std_logic_vector(92 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int93_t(x : std_logic_vector) return int93_t is
  variable rv : int93_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint94_t_to_slv(x : uint94_t) return std_logic_vector is
  variable rv : std_logic_vector(93 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint94_t(x : std_logic_vector) return uint94_t is
  variable rv : uint94_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int94_t_to_slv(x : int94_t) return std_logic_vector is
  variable rv : std_logic_vector(93 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int94_t(x : std_logic_vector) return int94_t is
  variable rv : int94_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint95_t_to_slv(x : uint95_t) return std_logic_vector is
  variable rv : std_logic_vector(94 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint95_t(x : std_logic_vector) return uint95_t is
  variable rv : uint95_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int95_t_to_slv(x : int95_t) return std_logic_vector is
  variable rv : std_logic_vector(94 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int95_t(x : std_logic_vector) return int95_t is
  variable rv : int95_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint96_t_to_slv(x : uint96_t) return std_logic_vector is
  variable rv : std_logic_vector(95 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint96_t(x : std_logic_vector) return uint96_t is
  variable rv : uint96_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int96_t_to_slv(x : int96_t) return std_logic_vector is
  variable rv : std_logic_vector(95 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int96_t(x : std_logic_vector) return int96_t is
  variable rv : int96_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint97_t_to_slv(x : uint97_t) return std_logic_vector is
  variable rv : std_logic_vector(96 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint97_t(x : std_logic_vector) return uint97_t is
  variable rv : uint97_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int97_t_to_slv(x : int97_t) return std_logic_vector is
  variable rv : std_logic_vector(96 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int97_t(x : std_logic_vector) return int97_t is
  variable rv : int97_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint98_t_to_slv(x : uint98_t) return std_logic_vector is
  variable rv : std_logic_vector(97 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint98_t(x : std_logic_vector) return uint98_t is
  variable rv : uint98_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int98_t_to_slv(x : int98_t) return std_logic_vector is
  variable rv : std_logic_vector(97 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int98_t(x : std_logic_vector) return int98_t is
  variable rv : int98_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint99_t_to_slv(x : uint99_t) return std_logic_vector is
  variable rv : std_logic_vector(98 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint99_t(x : std_logic_vector) return uint99_t is
  variable rv : uint99_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int99_t_to_slv(x : int99_t) return std_logic_vector is
  variable rv : std_logic_vector(98 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int99_t(x : std_logic_vector) return int99_t is
  variable rv : int99_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint100_t_to_slv(x : uint100_t) return std_logic_vector is
  variable rv : std_logic_vector(99 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint100_t(x : std_logic_vector) return uint100_t is
  variable rv : uint100_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int100_t_to_slv(x : int100_t) return std_logic_vector is
  variable rv : std_logic_vector(99 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int100_t(x : std_logic_vector) return int100_t is
  variable rv : int100_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint101_t_to_slv(x : uint101_t) return std_logic_vector is
  variable rv : std_logic_vector(100 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint101_t(x : std_logic_vector) return uint101_t is
  variable rv : uint101_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int101_t_to_slv(x : int101_t) return std_logic_vector is
  variable rv : std_logic_vector(100 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int101_t(x : std_logic_vector) return int101_t is
  variable rv : int101_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint102_t_to_slv(x : uint102_t) return std_logic_vector is
  variable rv : std_logic_vector(101 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint102_t(x : std_logic_vector) return uint102_t is
  variable rv : uint102_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int102_t_to_slv(x : int102_t) return std_logic_vector is
  variable rv : std_logic_vector(101 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int102_t(x : std_logic_vector) return int102_t is
  variable rv : int102_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint103_t_to_slv(x : uint103_t) return std_logic_vector is
  variable rv : std_logic_vector(102 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint103_t(x : std_logic_vector) return uint103_t is
  variable rv : uint103_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int103_t_to_slv(x : int103_t) return std_logic_vector is
  variable rv : std_logic_vector(102 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int103_t(x : std_logic_vector) return int103_t is
  variable rv : int103_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint104_t_to_slv(x : uint104_t) return std_logic_vector is
  variable rv : std_logic_vector(103 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint104_t(x : std_logic_vector) return uint104_t is
  variable rv : uint104_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int104_t_to_slv(x : int104_t) return std_logic_vector is
  variable rv : std_logic_vector(103 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int104_t(x : std_logic_vector) return int104_t is
  variable rv : int104_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint105_t_to_slv(x : uint105_t) return std_logic_vector is
  variable rv : std_logic_vector(104 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint105_t(x : std_logic_vector) return uint105_t is
  variable rv : uint105_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int105_t_to_slv(x : int105_t) return std_logic_vector is
  variable rv : std_logic_vector(104 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int105_t(x : std_logic_vector) return int105_t is
  variable rv : int105_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint106_t_to_slv(x : uint106_t) return std_logic_vector is
  variable rv : std_logic_vector(105 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint106_t(x : std_logic_vector) return uint106_t is
  variable rv : uint106_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int106_t_to_slv(x : int106_t) return std_logic_vector is
  variable rv : std_logic_vector(105 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int106_t(x : std_logic_vector) return int106_t is
  variable rv : int106_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint107_t_to_slv(x : uint107_t) return std_logic_vector is
  variable rv : std_logic_vector(106 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint107_t(x : std_logic_vector) return uint107_t is
  variable rv : uint107_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int107_t_to_slv(x : int107_t) return std_logic_vector is
  variable rv : std_logic_vector(106 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int107_t(x : std_logic_vector) return int107_t is
  variable rv : int107_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint108_t_to_slv(x : uint108_t) return std_logic_vector is
  variable rv : std_logic_vector(107 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint108_t(x : std_logic_vector) return uint108_t is
  variable rv : uint108_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int108_t_to_slv(x : int108_t) return std_logic_vector is
  variable rv : std_logic_vector(107 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int108_t(x : std_logic_vector) return int108_t is
  variable rv : int108_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint109_t_to_slv(x : uint109_t) return std_logic_vector is
  variable rv : std_logic_vector(108 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint109_t(x : std_logic_vector) return uint109_t is
  variable rv : uint109_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int109_t_to_slv(x : int109_t) return std_logic_vector is
  variable rv : std_logic_vector(108 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int109_t(x : std_logic_vector) return int109_t is
  variable rv : int109_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint110_t_to_slv(x : uint110_t) return std_logic_vector is
  variable rv : std_logic_vector(109 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint110_t(x : std_logic_vector) return uint110_t is
  variable rv : uint110_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int110_t_to_slv(x : int110_t) return std_logic_vector is
  variable rv : std_logic_vector(109 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int110_t(x : std_logic_vector) return int110_t is
  variable rv : int110_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint111_t_to_slv(x : uint111_t) return std_logic_vector is
  variable rv : std_logic_vector(110 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint111_t(x : std_logic_vector) return uint111_t is
  variable rv : uint111_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int111_t_to_slv(x : int111_t) return std_logic_vector is
  variable rv : std_logic_vector(110 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int111_t(x : std_logic_vector) return int111_t is
  variable rv : int111_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint112_t_to_slv(x : uint112_t) return std_logic_vector is
  variable rv : std_logic_vector(111 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint112_t(x : std_logic_vector) return uint112_t is
  variable rv : uint112_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int112_t_to_slv(x : int112_t) return std_logic_vector is
  variable rv : std_logic_vector(111 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int112_t(x : std_logic_vector) return int112_t is
  variable rv : int112_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint113_t_to_slv(x : uint113_t) return std_logic_vector is
  variable rv : std_logic_vector(112 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint113_t(x : std_logic_vector) return uint113_t is
  variable rv : uint113_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int113_t_to_slv(x : int113_t) return std_logic_vector is
  variable rv : std_logic_vector(112 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int113_t(x : std_logic_vector) return int113_t is
  variable rv : int113_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint114_t_to_slv(x : uint114_t) return std_logic_vector is
  variable rv : std_logic_vector(113 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint114_t(x : std_logic_vector) return uint114_t is
  variable rv : uint114_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int114_t_to_slv(x : int114_t) return std_logic_vector is
  variable rv : std_logic_vector(113 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int114_t(x : std_logic_vector) return int114_t is
  variable rv : int114_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint115_t_to_slv(x : uint115_t) return std_logic_vector is
  variable rv : std_logic_vector(114 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint115_t(x : std_logic_vector) return uint115_t is
  variable rv : uint115_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int115_t_to_slv(x : int115_t) return std_logic_vector is
  variable rv : std_logic_vector(114 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int115_t(x : std_logic_vector) return int115_t is
  variable rv : int115_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint116_t_to_slv(x : uint116_t) return std_logic_vector is
  variable rv : std_logic_vector(115 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint116_t(x : std_logic_vector) return uint116_t is
  variable rv : uint116_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int116_t_to_slv(x : int116_t) return std_logic_vector is
  variable rv : std_logic_vector(115 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int116_t(x : std_logic_vector) return int116_t is
  variable rv : int116_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint117_t_to_slv(x : uint117_t) return std_logic_vector is
  variable rv : std_logic_vector(116 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint117_t(x : std_logic_vector) return uint117_t is
  variable rv : uint117_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int117_t_to_slv(x : int117_t) return std_logic_vector is
  variable rv : std_logic_vector(116 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int117_t(x : std_logic_vector) return int117_t is
  variable rv : int117_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint118_t_to_slv(x : uint118_t) return std_logic_vector is
  variable rv : std_logic_vector(117 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint118_t(x : std_logic_vector) return uint118_t is
  variable rv : uint118_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int118_t_to_slv(x : int118_t) return std_logic_vector is
  variable rv : std_logic_vector(117 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int118_t(x : std_logic_vector) return int118_t is
  variable rv : int118_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint119_t_to_slv(x : uint119_t) return std_logic_vector is
  variable rv : std_logic_vector(118 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint119_t(x : std_logic_vector) return uint119_t is
  variable rv : uint119_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int119_t_to_slv(x : int119_t) return std_logic_vector is
  variable rv : std_logic_vector(118 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int119_t(x : std_logic_vector) return int119_t is
  variable rv : int119_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint120_t_to_slv(x : uint120_t) return std_logic_vector is
  variable rv : std_logic_vector(119 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint120_t(x : std_logic_vector) return uint120_t is
  variable rv : uint120_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int120_t_to_slv(x : int120_t) return std_logic_vector is
  variable rv : std_logic_vector(119 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int120_t(x : std_logic_vector) return int120_t is
  variable rv : int120_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint121_t_to_slv(x : uint121_t) return std_logic_vector is
  variable rv : std_logic_vector(120 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint121_t(x : std_logic_vector) return uint121_t is
  variable rv : uint121_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int121_t_to_slv(x : int121_t) return std_logic_vector is
  variable rv : std_logic_vector(120 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int121_t(x : std_logic_vector) return int121_t is
  variable rv : int121_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint122_t_to_slv(x : uint122_t) return std_logic_vector is
  variable rv : std_logic_vector(121 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint122_t(x : std_logic_vector) return uint122_t is
  variable rv : uint122_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int122_t_to_slv(x : int122_t) return std_logic_vector is
  variable rv : std_logic_vector(121 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int122_t(x : std_logic_vector) return int122_t is
  variable rv : int122_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint123_t_to_slv(x : uint123_t) return std_logic_vector is
  variable rv : std_logic_vector(122 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint123_t(x : std_logic_vector) return uint123_t is
  variable rv : uint123_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int123_t_to_slv(x : int123_t) return std_logic_vector is
  variable rv : std_logic_vector(122 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int123_t(x : std_logic_vector) return int123_t is
  variable rv : int123_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint124_t_to_slv(x : uint124_t) return std_logic_vector is
  variable rv : std_logic_vector(123 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint124_t(x : std_logic_vector) return uint124_t is
  variable rv : uint124_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int124_t_to_slv(x : int124_t) return std_logic_vector is
  variable rv : std_logic_vector(123 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int124_t(x : std_logic_vector) return int124_t is
  variable rv : int124_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint125_t_to_slv(x : uint125_t) return std_logic_vector is
  variable rv : std_logic_vector(124 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint125_t(x : std_logic_vector) return uint125_t is
  variable rv : uint125_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int125_t_to_slv(x : int125_t) return std_logic_vector is
  variable rv : std_logic_vector(124 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int125_t(x : std_logic_vector) return int125_t is
  variable rv : int125_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint126_t_to_slv(x : uint126_t) return std_logic_vector is
  variable rv : std_logic_vector(125 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint126_t(x : std_logic_vector) return uint126_t is
  variable rv : uint126_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int126_t_to_slv(x : int126_t) return std_logic_vector is
  variable rv : std_logic_vector(125 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int126_t(x : std_logic_vector) return int126_t is
  variable rv : int126_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint127_t_to_slv(x : uint127_t) return std_logic_vector is
  variable rv : std_logic_vector(126 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint127_t(x : std_logic_vector) return uint127_t is
  variable rv : uint127_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int127_t_to_slv(x : int127_t) return std_logic_vector is
  variable rv : std_logic_vector(126 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int127_t(x : std_logic_vector) return int127_t is
  variable rv : int127_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint128_t_to_slv(x : uint128_t) return std_logic_vector is
  variable rv : std_logic_vector(127 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint128_t(x : std_logic_vector) return uint128_t is
  variable rv : uint128_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int128_t_to_slv(x : int128_t) return std_logic_vector is
  variable rv : std_logic_vector(127 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int128_t(x : std_logic_vector) return int128_t is
  variable rv : int128_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint129_t_to_slv(x : uint129_t) return std_logic_vector is
  variable rv : std_logic_vector(128 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint129_t(x : std_logic_vector) return uint129_t is
  variable rv : uint129_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int129_t_to_slv(x : int129_t) return std_logic_vector is
  variable rv : std_logic_vector(128 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int129_t(x : std_logic_vector) return int129_t is
  variable rv : int129_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint130_t_to_slv(x : uint130_t) return std_logic_vector is
  variable rv : std_logic_vector(129 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint130_t(x : std_logic_vector) return uint130_t is
  variable rv : uint130_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int130_t_to_slv(x : int130_t) return std_logic_vector is
  variable rv : std_logic_vector(129 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int130_t(x : std_logic_vector) return int130_t is
  variable rv : int130_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint131_t_to_slv(x : uint131_t) return std_logic_vector is
  variable rv : std_logic_vector(130 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint131_t(x : std_logic_vector) return uint131_t is
  variable rv : uint131_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int131_t_to_slv(x : int131_t) return std_logic_vector is
  variable rv : std_logic_vector(130 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int131_t(x : std_logic_vector) return int131_t is
  variable rv : int131_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint132_t_to_slv(x : uint132_t) return std_logic_vector is
  variable rv : std_logic_vector(131 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint132_t(x : std_logic_vector) return uint132_t is
  variable rv : uint132_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int132_t_to_slv(x : int132_t) return std_logic_vector is
  variable rv : std_logic_vector(131 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int132_t(x : std_logic_vector) return int132_t is
  variable rv : int132_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint133_t_to_slv(x : uint133_t) return std_logic_vector is
  variable rv : std_logic_vector(132 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint133_t(x : std_logic_vector) return uint133_t is
  variable rv : uint133_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int133_t_to_slv(x : int133_t) return std_logic_vector is
  variable rv : std_logic_vector(132 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int133_t(x : std_logic_vector) return int133_t is
  variable rv : int133_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint134_t_to_slv(x : uint134_t) return std_logic_vector is
  variable rv : std_logic_vector(133 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint134_t(x : std_logic_vector) return uint134_t is
  variable rv : uint134_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int134_t_to_slv(x : int134_t) return std_logic_vector is
  variable rv : std_logic_vector(133 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int134_t(x : std_logic_vector) return int134_t is
  variable rv : int134_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint135_t_to_slv(x : uint135_t) return std_logic_vector is
  variable rv : std_logic_vector(134 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint135_t(x : std_logic_vector) return uint135_t is
  variable rv : uint135_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int135_t_to_slv(x : int135_t) return std_logic_vector is
  variable rv : std_logic_vector(134 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int135_t(x : std_logic_vector) return int135_t is
  variable rv : int135_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint136_t_to_slv(x : uint136_t) return std_logic_vector is
  variable rv : std_logic_vector(135 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint136_t(x : std_logic_vector) return uint136_t is
  variable rv : uint136_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int136_t_to_slv(x : int136_t) return std_logic_vector is
  variable rv : std_logic_vector(135 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int136_t(x : std_logic_vector) return int136_t is
  variable rv : int136_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint137_t_to_slv(x : uint137_t) return std_logic_vector is
  variable rv : std_logic_vector(136 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint137_t(x : std_logic_vector) return uint137_t is
  variable rv : uint137_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int137_t_to_slv(x : int137_t) return std_logic_vector is
  variable rv : std_logic_vector(136 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int137_t(x : std_logic_vector) return int137_t is
  variable rv : int137_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint138_t_to_slv(x : uint138_t) return std_logic_vector is
  variable rv : std_logic_vector(137 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint138_t(x : std_logic_vector) return uint138_t is
  variable rv : uint138_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int138_t_to_slv(x : int138_t) return std_logic_vector is
  variable rv : std_logic_vector(137 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int138_t(x : std_logic_vector) return int138_t is
  variable rv : int138_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint139_t_to_slv(x : uint139_t) return std_logic_vector is
  variable rv : std_logic_vector(138 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint139_t(x : std_logic_vector) return uint139_t is
  variable rv : uint139_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int139_t_to_slv(x : int139_t) return std_logic_vector is
  variable rv : std_logic_vector(138 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int139_t(x : std_logic_vector) return int139_t is
  variable rv : int139_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint140_t_to_slv(x : uint140_t) return std_logic_vector is
  variable rv : std_logic_vector(139 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint140_t(x : std_logic_vector) return uint140_t is
  variable rv : uint140_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int140_t_to_slv(x : int140_t) return std_logic_vector is
  variable rv : std_logic_vector(139 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int140_t(x : std_logic_vector) return int140_t is
  variable rv : int140_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint141_t_to_slv(x : uint141_t) return std_logic_vector is
  variable rv : std_logic_vector(140 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint141_t(x : std_logic_vector) return uint141_t is
  variable rv : uint141_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int141_t_to_slv(x : int141_t) return std_logic_vector is
  variable rv : std_logic_vector(140 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int141_t(x : std_logic_vector) return int141_t is
  variable rv : int141_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint142_t_to_slv(x : uint142_t) return std_logic_vector is
  variable rv : std_logic_vector(141 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint142_t(x : std_logic_vector) return uint142_t is
  variable rv : uint142_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int142_t_to_slv(x : int142_t) return std_logic_vector is
  variable rv : std_logic_vector(141 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int142_t(x : std_logic_vector) return int142_t is
  variable rv : int142_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint143_t_to_slv(x : uint143_t) return std_logic_vector is
  variable rv : std_logic_vector(142 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint143_t(x : std_logic_vector) return uint143_t is
  variable rv : uint143_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int143_t_to_slv(x : int143_t) return std_logic_vector is
  variable rv : std_logic_vector(142 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int143_t(x : std_logic_vector) return int143_t is
  variable rv : int143_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint144_t_to_slv(x : uint144_t) return std_logic_vector is
  variable rv : std_logic_vector(143 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint144_t(x : std_logic_vector) return uint144_t is
  variable rv : uint144_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int144_t_to_slv(x : int144_t) return std_logic_vector is
  variable rv : std_logic_vector(143 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int144_t(x : std_logic_vector) return int144_t is
  variable rv : int144_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint145_t_to_slv(x : uint145_t) return std_logic_vector is
  variable rv : std_logic_vector(144 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint145_t(x : std_logic_vector) return uint145_t is
  variable rv : uint145_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int145_t_to_slv(x : int145_t) return std_logic_vector is
  variable rv : std_logic_vector(144 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int145_t(x : std_logic_vector) return int145_t is
  variable rv : int145_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint146_t_to_slv(x : uint146_t) return std_logic_vector is
  variable rv : std_logic_vector(145 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint146_t(x : std_logic_vector) return uint146_t is
  variable rv : uint146_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int146_t_to_slv(x : int146_t) return std_logic_vector is
  variable rv : std_logic_vector(145 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int146_t(x : std_logic_vector) return int146_t is
  variable rv : int146_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint147_t_to_slv(x : uint147_t) return std_logic_vector is
  variable rv : std_logic_vector(146 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint147_t(x : std_logic_vector) return uint147_t is
  variable rv : uint147_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int147_t_to_slv(x : int147_t) return std_logic_vector is
  variable rv : std_logic_vector(146 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int147_t(x : std_logic_vector) return int147_t is
  variable rv : int147_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint148_t_to_slv(x : uint148_t) return std_logic_vector is
  variable rv : std_logic_vector(147 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint148_t(x : std_logic_vector) return uint148_t is
  variable rv : uint148_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int148_t_to_slv(x : int148_t) return std_logic_vector is
  variable rv : std_logic_vector(147 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int148_t(x : std_logic_vector) return int148_t is
  variable rv : int148_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint149_t_to_slv(x : uint149_t) return std_logic_vector is
  variable rv : std_logic_vector(148 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint149_t(x : std_logic_vector) return uint149_t is
  variable rv : uint149_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int149_t_to_slv(x : int149_t) return std_logic_vector is
  variable rv : std_logic_vector(148 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int149_t(x : std_logic_vector) return int149_t is
  variable rv : int149_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint150_t_to_slv(x : uint150_t) return std_logic_vector is
  variable rv : std_logic_vector(149 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint150_t(x : std_logic_vector) return uint150_t is
  variable rv : uint150_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int150_t_to_slv(x : int150_t) return std_logic_vector is
  variable rv : std_logic_vector(149 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int150_t(x : std_logic_vector) return int150_t is
  variable rv : int150_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint151_t_to_slv(x : uint151_t) return std_logic_vector is
  variable rv : std_logic_vector(150 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint151_t(x : std_logic_vector) return uint151_t is
  variable rv : uint151_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int151_t_to_slv(x : int151_t) return std_logic_vector is
  variable rv : std_logic_vector(150 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int151_t(x : std_logic_vector) return int151_t is
  variable rv : int151_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint152_t_to_slv(x : uint152_t) return std_logic_vector is
  variable rv : std_logic_vector(151 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint152_t(x : std_logic_vector) return uint152_t is
  variable rv : uint152_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int152_t_to_slv(x : int152_t) return std_logic_vector is
  variable rv : std_logic_vector(151 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int152_t(x : std_logic_vector) return int152_t is
  variable rv : int152_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint153_t_to_slv(x : uint153_t) return std_logic_vector is
  variable rv : std_logic_vector(152 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint153_t(x : std_logic_vector) return uint153_t is
  variable rv : uint153_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int153_t_to_slv(x : int153_t) return std_logic_vector is
  variable rv : std_logic_vector(152 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int153_t(x : std_logic_vector) return int153_t is
  variable rv : int153_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint154_t_to_slv(x : uint154_t) return std_logic_vector is
  variable rv : std_logic_vector(153 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint154_t(x : std_logic_vector) return uint154_t is
  variable rv : uint154_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int154_t_to_slv(x : int154_t) return std_logic_vector is
  variable rv : std_logic_vector(153 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int154_t(x : std_logic_vector) return int154_t is
  variable rv : int154_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint155_t_to_slv(x : uint155_t) return std_logic_vector is
  variable rv : std_logic_vector(154 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint155_t(x : std_logic_vector) return uint155_t is
  variable rv : uint155_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int155_t_to_slv(x : int155_t) return std_logic_vector is
  variable rv : std_logic_vector(154 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int155_t(x : std_logic_vector) return int155_t is
  variable rv : int155_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint156_t_to_slv(x : uint156_t) return std_logic_vector is
  variable rv : std_logic_vector(155 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint156_t(x : std_logic_vector) return uint156_t is
  variable rv : uint156_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int156_t_to_slv(x : int156_t) return std_logic_vector is
  variable rv : std_logic_vector(155 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int156_t(x : std_logic_vector) return int156_t is
  variable rv : int156_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint157_t_to_slv(x : uint157_t) return std_logic_vector is
  variable rv : std_logic_vector(156 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint157_t(x : std_logic_vector) return uint157_t is
  variable rv : uint157_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int157_t_to_slv(x : int157_t) return std_logic_vector is
  variable rv : std_logic_vector(156 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int157_t(x : std_logic_vector) return int157_t is
  variable rv : int157_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint158_t_to_slv(x : uint158_t) return std_logic_vector is
  variable rv : std_logic_vector(157 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint158_t(x : std_logic_vector) return uint158_t is
  variable rv : uint158_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int158_t_to_slv(x : int158_t) return std_logic_vector is
  variable rv : std_logic_vector(157 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int158_t(x : std_logic_vector) return int158_t is
  variable rv : int158_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint159_t_to_slv(x : uint159_t) return std_logic_vector is
  variable rv : std_logic_vector(158 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint159_t(x : std_logic_vector) return uint159_t is
  variable rv : uint159_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int159_t_to_slv(x : int159_t) return std_logic_vector is
  variable rv : std_logic_vector(158 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int159_t(x : std_logic_vector) return int159_t is
  variable rv : int159_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint160_t_to_slv(x : uint160_t) return std_logic_vector is
  variable rv : std_logic_vector(159 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint160_t(x : std_logic_vector) return uint160_t is
  variable rv : uint160_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int160_t_to_slv(x : int160_t) return std_logic_vector is
  variable rv : std_logic_vector(159 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int160_t(x : std_logic_vector) return int160_t is
  variable rv : int160_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint161_t_to_slv(x : uint161_t) return std_logic_vector is
  variable rv : std_logic_vector(160 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint161_t(x : std_logic_vector) return uint161_t is
  variable rv : uint161_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int161_t_to_slv(x : int161_t) return std_logic_vector is
  variable rv : std_logic_vector(160 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int161_t(x : std_logic_vector) return int161_t is
  variable rv : int161_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint162_t_to_slv(x : uint162_t) return std_logic_vector is
  variable rv : std_logic_vector(161 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint162_t(x : std_logic_vector) return uint162_t is
  variable rv : uint162_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int162_t_to_slv(x : int162_t) return std_logic_vector is
  variable rv : std_logic_vector(161 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int162_t(x : std_logic_vector) return int162_t is
  variable rv : int162_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint163_t_to_slv(x : uint163_t) return std_logic_vector is
  variable rv : std_logic_vector(162 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint163_t(x : std_logic_vector) return uint163_t is
  variable rv : uint163_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int163_t_to_slv(x : int163_t) return std_logic_vector is
  variable rv : std_logic_vector(162 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int163_t(x : std_logic_vector) return int163_t is
  variable rv : int163_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint164_t_to_slv(x : uint164_t) return std_logic_vector is
  variable rv : std_logic_vector(163 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint164_t(x : std_logic_vector) return uint164_t is
  variable rv : uint164_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int164_t_to_slv(x : int164_t) return std_logic_vector is
  variable rv : std_logic_vector(163 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int164_t(x : std_logic_vector) return int164_t is
  variable rv : int164_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint165_t_to_slv(x : uint165_t) return std_logic_vector is
  variable rv : std_logic_vector(164 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint165_t(x : std_logic_vector) return uint165_t is
  variable rv : uint165_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int165_t_to_slv(x : int165_t) return std_logic_vector is
  variable rv : std_logic_vector(164 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int165_t(x : std_logic_vector) return int165_t is
  variable rv : int165_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint166_t_to_slv(x : uint166_t) return std_logic_vector is
  variable rv : std_logic_vector(165 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint166_t(x : std_logic_vector) return uint166_t is
  variable rv : uint166_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int166_t_to_slv(x : int166_t) return std_logic_vector is
  variable rv : std_logic_vector(165 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int166_t(x : std_logic_vector) return int166_t is
  variable rv : int166_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint167_t_to_slv(x : uint167_t) return std_logic_vector is
  variable rv : std_logic_vector(166 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint167_t(x : std_logic_vector) return uint167_t is
  variable rv : uint167_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int167_t_to_slv(x : int167_t) return std_logic_vector is
  variable rv : std_logic_vector(166 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int167_t(x : std_logic_vector) return int167_t is
  variable rv : int167_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint168_t_to_slv(x : uint168_t) return std_logic_vector is
  variable rv : std_logic_vector(167 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint168_t(x : std_logic_vector) return uint168_t is
  variable rv : uint168_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int168_t_to_slv(x : int168_t) return std_logic_vector is
  variable rv : std_logic_vector(167 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int168_t(x : std_logic_vector) return int168_t is
  variable rv : int168_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint169_t_to_slv(x : uint169_t) return std_logic_vector is
  variable rv : std_logic_vector(168 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint169_t(x : std_logic_vector) return uint169_t is
  variable rv : uint169_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int169_t_to_slv(x : int169_t) return std_logic_vector is
  variable rv : std_logic_vector(168 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int169_t(x : std_logic_vector) return int169_t is
  variable rv : int169_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint170_t_to_slv(x : uint170_t) return std_logic_vector is
  variable rv : std_logic_vector(169 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint170_t(x : std_logic_vector) return uint170_t is
  variable rv : uint170_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int170_t_to_slv(x : int170_t) return std_logic_vector is
  variable rv : std_logic_vector(169 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int170_t(x : std_logic_vector) return int170_t is
  variable rv : int170_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint171_t_to_slv(x : uint171_t) return std_logic_vector is
  variable rv : std_logic_vector(170 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint171_t(x : std_logic_vector) return uint171_t is
  variable rv : uint171_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int171_t_to_slv(x : int171_t) return std_logic_vector is
  variable rv : std_logic_vector(170 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int171_t(x : std_logic_vector) return int171_t is
  variable rv : int171_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint172_t_to_slv(x : uint172_t) return std_logic_vector is
  variable rv : std_logic_vector(171 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint172_t(x : std_logic_vector) return uint172_t is
  variable rv : uint172_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int172_t_to_slv(x : int172_t) return std_logic_vector is
  variable rv : std_logic_vector(171 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int172_t(x : std_logic_vector) return int172_t is
  variable rv : int172_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint173_t_to_slv(x : uint173_t) return std_logic_vector is
  variable rv : std_logic_vector(172 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint173_t(x : std_logic_vector) return uint173_t is
  variable rv : uint173_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int173_t_to_slv(x : int173_t) return std_logic_vector is
  variable rv : std_logic_vector(172 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int173_t(x : std_logic_vector) return int173_t is
  variable rv : int173_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint174_t_to_slv(x : uint174_t) return std_logic_vector is
  variable rv : std_logic_vector(173 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint174_t(x : std_logic_vector) return uint174_t is
  variable rv : uint174_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int174_t_to_slv(x : int174_t) return std_logic_vector is
  variable rv : std_logic_vector(173 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int174_t(x : std_logic_vector) return int174_t is
  variable rv : int174_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint175_t_to_slv(x : uint175_t) return std_logic_vector is
  variable rv : std_logic_vector(174 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint175_t(x : std_logic_vector) return uint175_t is
  variable rv : uint175_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int175_t_to_slv(x : int175_t) return std_logic_vector is
  variable rv : std_logic_vector(174 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int175_t(x : std_logic_vector) return int175_t is
  variable rv : int175_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint176_t_to_slv(x : uint176_t) return std_logic_vector is
  variable rv : std_logic_vector(175 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint176_t(x : std_logic_vector) return uint176_t is
  variable rv : uint176_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int176_t_to_slv(x : int176_t) return std_logic_vector is
  variable rv : std_logic_vector(175 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int176_t(x : std_logic_vector) return int176_t is
  variable rv : int176_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint177_t_to_slv(x : uint177_t) return std_logic_vector is
  variable rv : std_logic_vector(176 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint177_t(x : std_logic_vector) return uint177_t is
  variable rv : uint177_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int177_t_to_slv(x : int177_t) return std_logic_vector is
  variable rv : std_logic_vector(176 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int177_t(x : std_logic_vector) return int177_t is
  variable rv : int177_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint178_t_to_slv(x : uint178_t) return std_logic_vector is
  variable rv : std_logic_vector(177 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint178_t(x : std_logic_vector) return uint178_t is
  variable rv : uint178_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int178_t_to_slv(x : int178_t) return std_logic_vector is
  variable rv : std_logic_vector(177 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int178_t(x : std_logic_vector) return int178_t is
  variable rv : int178_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint179_t_to_slv(x : uint179_t) return std_logic_vector is
  variable rv : std_logic_vector(178 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint179_t(x : std_logic_vector) return uint179_t is
  variable rv : uint179_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int179_t_to_slv(x : int179_t) return std_logic_vector is
  variable rv : std_logic_vector(178 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int179_t(x : std_logic_vector) return int179_t is
  variable rv : int179_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint180_t_to_slv(x : uint180_t) return std_logic_vector is
  variable rv : std_logic_vector(179 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint180_t(x : std_logic_vector) return uint180_t is
  variable rv : uint180_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int180_t_to_slv(x : int180_t) return std_logic_vector is
  variable rv : std_logic_vector(179 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int180_t(x : std_logic_vector) return int180_t is
  variable rv : int180_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint181_t_to_slv(x : uint181_t) return std_logic_vector is
  variable rv : std_logic_vector(180 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint181_t(x : std_logic_vector) return uint181_t is
  variable rv : uint181_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int181_t_to_slv(x : int181_t) return std_logic_vector is
  variable rv : std_logic_vector(180 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int181_t(x : std_logic_vector) return int181_t is
  variable rv : int181_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint182_t_to_slv(x : uint182_t) return std_logic_vector is
  variable rv : std_logic_vector(181 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint182_t(x : std_logic_vector) return uint182_t is
  variable rv : uint182_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int182_t_to_slv(x : int182_t) return std_logic_vector is
  variable rv : std_logic_vector(181 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int182_t(x : std_logic_vector) return int182_t is
  variable rv : int182_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint183_t_to_slv(x : uint183_t) return std_logic_vector is
  variable rv : std_logic_vector(182 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint183_t(x : std_logic_vector) return uint183_t is
  variable rv : uint183_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int183_t_to_slv(x : int183_t) return std_logic_vector is
  variable rv : std_logic_vector(182 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int183_t(x : std_logic_vector) return int183_t is
  variable rv : int183_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint184_t_to_slv(x : uint184_t) return std_logic_vector is
  variable rv : std_logic_vector(183 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint184_t(x : std_logic_vector) return uint184_t is
  variable rv : uint184_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int184_t_to_slv(x : int184_t) return std_logic_vector is
  variable rv : std_logic_vector(183 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int184_t(x : std_logic_vector) return int184_t is
  variable rv : int184_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint185_t_to_slv(x : uint185_t) return std_logic_vector is
  variable rv : std_logic_vector(184 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint185_t(x : std_logic_vector) return uint185_t is
  variable rv : uint185_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int185_t_to_slv(x : int185_t) return std_logic_vector is
  variable rv : std_logic_vector(184 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int185_t(x : std_logic_vector) return int185_t is
  variable rv : int185_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint186_t_to_slv(x : uint186_t) return std_logic_vector is
  variable rv : std_logic_vector(185 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint186_t(x : std_logic_vector) return uint186_t is
  variable rv : uint186_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int186_t_to_slv(x : int186_t) return std_logic_vector is
  variable rv : std_logic_vector(185 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int186_t(x : std_logic_vector) return int186_t is
  variable rv : int186_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint187_t_to_slv(x : uint187_t) return std_logic_vector is
  variable rv : std_logic_vector(186 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint187_t(x : std_logic_vector) return uint187_t is
  variable rv : uint187_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int187_t_to_slv(x : int187_t) return std_logic_vector is
  variable rv : std_logic_vector(186 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int187_t(x : std_logic_vector) return int187_t is
  variable rv : int187_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint188_t_to_slv(x : uint188_t) return std_logic_vector is
  variable rv : std_logic_vector(187 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint188_t(x : std_logic_vector) return uint188_t is
  variable rv : uint188_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int188_t_to_slv(x : int188_t) return std_logic_vector is
  variable rv : std_logic_vector(187 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int188_t(x : std_logic_vector) return int188_t is
  variable rv : int188_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint189_t_to_slv(x : uint189_t) return std_logic_vector is
  variable rv : std_logic_vector(188 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint189_t(x : std_logic_vector) return uint189_t is
  variable rv : uint189_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int189_t_to_slv(x : int189_t) return std_logic_vector is
  variable rv : std_logic_vector(188 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int189_t(x : std_logic_vector) return int189_t is
  variable rv : int189_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint190_t_to_slv(x : uint190_t) return std_logic_vector is
  variable rv : std_logic_vector(189 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint190_t(x : std_logic_vector) return uint190_t is
  variable rv : uint190_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int190_t_to_slv(x : int190_t) return std_logic_vector is
  variable rv : std_logic_vector(189 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int190_t(x : std_logic_vector) return int190_t is
  variable rv : int190_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint191_t_to_slv(x : uint191_t) return std_logic_vector is
  variable rv : std_logic_vector(190 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint191_t(x : std_logic_vector) return uint191_t is
  variable rv : uint191_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int191_t_to_slv(x : int191_t) return std_logic_vector is
  variable rv : std_logic_vector(190 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int191_t(x : std_logic_vector) return int191_t is
  variable rv : int191_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint192_t_to_slv(x : uint192_t) return std_logic_vector is
  variable rv : std_logic_vector(191 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint192_t(x : std_logic_vector) return uint192_t is
  variable rv : uint192_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int192_t_to_slv(x : int192_t) return std_logic_vector is
  variable rv : std_logic_vector(191 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int192_t(x : std_logic_vector) return int192_t is
  variable rv : int192_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint193_t_to_slv(x : uint193_t) return std_logic_vector is
  variable rv : std_logic_vector(192 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint193_t(x : std_logic_vector) return uint193_t is
  variable rv : uint193_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int193_t_to_slv(x : int193_t) return std_logic_vector is
  variable rv : std_logic_vector(192 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int193_t(x : std_logic_vector) return int193_t is
  variable rv : int193_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint194_t_to_slv(x : uint194_t) return std_logic_vector is
  variable rv : std_logic_vector(193 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint194_t(x : std_logic_vector) return uint194_t is
  variable rv : uint194_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int194_t_to_slv(x : int194_t) return std_logic_vector is
  variable rv : std_logic_vector(193 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int194_t(x : std_logic_vector) return int194_t is
  variable rv : int194_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint195_t_to_slv(x : uint195_t) return std_logic_vector is
  variable rv : std_logic_vector(194 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint195_t(x : std_logic_vector) return uint195_t is
  variable rv : uint195_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int195_t_to_slv(x : int195_t) return std_logic_vector is
  variable rv : std_logic_vector(194 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int195_t(x : std_logic_vector) return int195_t is
  variable rv : int195_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint196_t_to_slv(x : uint196_t) return std_logic_vector is
  variable rv : std_logic_vector(195 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint196_t(x : std_logic_vector) return uint196_t is
  variable rv : uint196_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int196_t_to_slv(x : int196_t) return std_logic_vector is
  variable rv : std_logic_vector(195 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int196_t(x : std_logic_vector) return int196_t is
  variable rv : int196_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint197_t_to_slv(x : uint197_t) return std_logic_vector is
  variable rv : std_logic_vector(196 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint197_t(x : std_logic_vector) return uint197_t is
  variable rv : uint197_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int197_t_to_slv(x : int197_t) return std_logic_vector is
  variable rv : std_logic_vector(196 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int197_t(x : std_logic_vector) return int197_t is
  variable rv : int197_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint198_t_to_slv(x : uint198_t) return std_logic_vector is
  variable rv : std_logic_vector(197 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint198_t(x : std_logic_vector) return uint198_t is
  variable rv : uint198_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int198_t_to_slv(x : int198_t) return std_logic_vector is
  variable rv : std_logic_vector(197 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int198_t(x : std_logic_vector) return int198_t is
  variable rv : int198_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint199_t_to_slv(x : uint199_t) return std_logic_vector is
  variable rv : std_logic_vector(198 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint199_t(x : std_logic_vector) return uint199_t is
  variable rv : uint199_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int199_t_to_slv(x : int199_t) return std_logic_vector is
  variable rv : std_logic_vector(198 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int199_t(x : std_logic_vector) return int199_t is
  variable rv : int199_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint200_t_to_slv(x : uint200_t) return std_logic_vector is
  variable rv : std_logic_vector(199 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint200_t(x : std_logic_vector) return uint200_t is
  variable rv : uint200_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int200_t_to_slv(x : int200_t) return std_logic_vector is
  variable rv : std_logic_vector(199 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int200_t(x : std_logic_vector) return int200_t is
  variable rv : int200_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint201_t_to_slv(x : uint201_t) return std_logic_vector is
  variable rv : std_logic_vector(200 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint201_t(x : std_logic_vector) return uint201_t is
  variable rv : uint201_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int201_t_to_slv(x : int201_t) return std_logic_vector is
  variable rv : std_logic_vector(200 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int201_t(x : std_logic_vector) return int201_t is
  variable rv : int201_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint202_t_to_slv(x : uint202_t) return std_logic_vector is
  variable rv : std_logic_vector(201 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint202_t(x : std_logic_vector) return uint202_t is
  variable rv : uint202_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int202_t_to_slv(x : int202_t) return std_logic_vector is
  variable rv : std_logic_vector(201 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int202_t(x : std_logic_vector) return int202_t is
  variable rv : int202_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint203_t_to_slv(x : uint203_t) return std_logic_vector is
  variable rv : std_logic_vector(202 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint203_t(x : std_logic_vector) return uint203_t is
  variable rv : uint203_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int203_t_to_slv(x : int203_t) return std_logic_vector is
  variable rv : std_logic_vector(202 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int203_t(x : std_logic_vector) return int203_t is
  variable rv : int203_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint204_t_to_slv(x : uint204_t) return std_logic_vector is
  variable rv : std_logic_vector(203 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint204_t(x : std_logic_vector) return uint204_t is
  variable rv : uint204_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int204_t_to_slv(x : int204_t) return std_logic_vector is
  variable rv : std_logic_vector(203 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int204_t(x : std_logic_vector) return int204_t is
  variable rv : int204_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint205_t_to_slv(x : uint205_t) return std_logic_vector is
  variable rv : std_logic_vector(204 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint205_t(x : std_logic_vector) return uint205_t is
  variable rv : uint205_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int205_t_to_slv(x : int205_t) return std_logic_vector is
  variable rv : std_logic_vector(204 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int205_t(x : std_logic_vector) return int205_t is
  variable rv : int205_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint206_t_to_slv(x : uint206_t) return std_logic_vector is
  variable rv : std_logic_vector(205 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint206_t(x : std_logic_vector) return uint206_t is
  variable rv : uint206_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int206_t_to_slv(x : int206_t) return std_logic_vector is
  variable rv : std_logic_vector(205 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int206_t(x : std_logic_vector) return int206_t is
  variable rv : int206_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint207_t_to_slv(x : uint207_t) return std_logic_vector is
  variable rv : std_logic_vector(206 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint207_t(x : std_logic_vector) return uint207_t is
  variable rv : uint207_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int207_t_to_slv(x : int207_t) return std_logic_vector is
  variable rv : std_logic_vector(206 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int207_t(x : std_logic_vector) return int207_t is
  variable rv : int207_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint208_t_to_slv(x : uint208_t) return std_logic_vector is
  variable rv : std_logic_vector(207 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint208_t(x : std_logic_vector) return uint208_t is
  variable rv : uint208_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int208_t_to_slv(x : int208_t) return std_logic_vector is
  variable rv : std_logic_vector(207 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int208_t(x : std_logic_vector) return int208_t is
  variable rv : int208_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint209_t_to_slv(x : uint209_t) return std_logic_vector is
  variable rv : std_logic_vector(208 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint209_t(x : std_logic_vector) return uint209_t is
  variable rv : uint209_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int209_t_to_slv(x : int209_t) return std_logic_vector is
  variable rv : std_logic_vector(208 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int209_t(x : std_logic_vector) return int209_t is
  variable rv : int209_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint210_t_to_slv(x : uint210_t) return std_logic_vector is
  variable rv : std_logic_vector(209 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint210_t(x : std_logic_vector) return uint210_t is
  variable rv : uint210_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int210_t_to_slv(x : int210_t) return std_logic_vector is
  variable rv : std_logic_vector(209 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int210_t(x : std_logic_vector) return int210_t is
  variable rv : int210_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint211_t_to_slv(x : uint211_t) return std_logic_vector is
  variable rv : std_logic_vector(210 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint211_t(x : std_logic_vector) return uint211_t is
  variable rv : uint211_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int211_t_to_slv(x : int211_t) return std_logic_vector is
  variable rv : std_logic_vector(210 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int211_t(x : std_logic_vector) return int211_t is
  variable rv : int211_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint212_t_to_slv(x : uint212_t) return std_logic_vector is
  variable rv : std_logic_vector(211 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint212_t(x : std_logic_vector) return uint212_t is
  variable rv : uint212_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int212_t_to_slv(x : int212_t) return std_logic_vector is
  variable rv : std_logic_vector(211 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int212_t(x : std_logic_vector) return int212_t is
  variable rv : int212_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint213_t_to_slv(x : uint213_t) return std_logic_vector is
  variable rv : std_logic_vector(212 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint213_t(x : std_logic_vector) return uint213_t is
  variable rv : uint213_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int213_t_to_slv(x : int213_t) return std_logic_vector is
  variable rv : std_logic_vector(212 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int213_t(x : std_logic_vector) return int213_t is
  variable rv : int213_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint214_t_to_slv(x : uint214_t) return std_logic_vector is
  variable rv : std_logic_vector(213 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint214_t(x : std_logic_vector) return uint214_t is
  variable rv : uint214_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int214_t_to_slv(x : int214_t) return std_logic_vector is
  variable rv : std_logic_vector(213 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int214_t(x : std_logic_vector) return int214_t is
  variable rv : int214_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint215_t_to_slv(x : uint215_t) return std_logic_vector is
  variable rv : std_logic_vector(214 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint215_t(x : std_logic_vector) return uint215_t is
  variable rv : uint215_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int215_t_to_slv(x : int215_t) return std_logic_vector is
  variable rv : std_logic_vector(214 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int215_t(x : std_logic_vector) return int215_t is
  variable rv : int215_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint216_t_to_slv(x : uint216_t) return std_logic_vector is
  variable rv : std_logic_vector(215 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint216_t(x : std_logic_vector) return uint216_t is
  variable rv : uint216_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int216_t_to_slv(x : int216_t) return std_logic_vector is
  variable rv : std_logic_vector(215 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int216_t(x : std_logic_vector) return int216_t is
  variable rv : int216_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint217_t_to_slv(x : uint217_t) return std_logic_vector is
  variable rv : std_logic_vector(216 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint217_t(x : std_logic_vector) return uint217_t is
  variable rv : uint217_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int217_t_to_slv(x : int217_t) return std_logic_vector is
  variable rv : std_logic_vector(216 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int217_t(x : std_logic_vector) return int217_t is
  variable rv : int217_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint218_t_to_slv(x : uint218_t) return std_logic_vector is
  variable rv : std_logic_vector(217 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint218_t(x : std_logic_vector) return uint218_t is
  variable rv : uint218_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int218_t_to_slv(x : int218_t) return std_logic_vector is
  variable rv : std_logic_vector(217 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int218_t(x : std_logic_vector) return int218_t is
  variable rv : int218_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint219_t_to_slv(x : uint219_t) return std_logic_vector is
  variable rv : std_logic_vector(218 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint219_t(x : std_logic_vector) return uint219_t is
  variable rv : uint219_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int219_t_to_slv(x : int219_t) return std_logic_vector is
  variable rv : std_logic_vector(218 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int219_t(x : std_logic_vector) return int219_t is
  variable rv : int219_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint220_t_to_slv(x : uint220_t) return std_logic_vector is
  variable rv : std_logic_vector(219 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint220_t(x : std_logic_vector) return uint220_t is
  variable rv : uint220_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int220_t_to_slv(x : int220_t) return std_logic_vector is
  variable rv : std_logic_vector(219 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int220_t(x : std_logic_vector) return int220_t is
  variable rv : int220_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint221_t_to_slv(x : uint221_t) return std_logic_vector is
  variable rv : std_logic_vector(220 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint221_t(x : std_logic_vector) return uint221_t is
  variable rv : uint221_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int221_t_to_slv(x : int221_t) return std_logic_vector is
  variable rv : std_logic_vector(220 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int221_t(x : std_logic_vector) return int221_t is
  variable rv : int221_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint222_t_to_slv(x : uint222_t) return std_logic_vector is
  variable rv : std_logic_vector(221 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint222_t(x : std_logic_vector) return uint222_t is
  variable rv : uint222_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int222_t_to_slv(x : int222_t) return std_logic_vector is
  variable rv : std_logic_vector(221 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int222_t(x : std_logic_vector) return int222_t is
  variable rv : int222_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint223_t_to_slv(x : uint223_t) return std_logic_vector is
  variable rv : std_logic_vector(222 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint223_t(x : std_logic_vector) return uint223_t is
  variable rv : uint223_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int223_t_to_slv(x : int223_t) return std_logic_vector is
  variable rv : std_logic_vector(222 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int223_t(x : std_logic_vector) return int223_t is
  variable rv : int223_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint224_t_to_slv(x : uint224_t) return std_logic_vector is
  variable rv : std_logic_vector(223 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint224_t(x : std_logic_vector) return uint224_t is
  variable rv : uint224_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int224_t_to_slv(x : int224_t) return std_logic_vector is
  variable rv : std_logic_vector(223 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int224_t(x : std_logic_vector) return int224_t is
  variable rv : int224_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint225_t_to_slv(x : uint225_t) return std_logic_vector is
  variable rv : std_logic_vector(224 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint225_t(x : std_logic_vector) return uint225_t is
  variable rv : uint225_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int225_t_to_slv(x : int225_t) return std_logic_vector is
  variable rv : std_logic_vector(224 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int225_t(x : std_logic_vector) return int225_t is
  variable rv : int225_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint226_t_to_slv(x : uint226_t) return std_logic_vector is
  variable rv : std_logic_vector(225 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint226_t(x : std_logic_vector) return uint226_t is
  variable rv : uint226_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int226_t_to_slv(x : int226_t) return std_logic_vector is
  variable rv : std_logic_vector(225 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int226_t(x : std_logic_vector) return int226_t is
  variable rv : int226_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint227_t_to_slv(x : uint227_t) return std_logic_vector is
  variable rv : std_logic_vector(226 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint227_t(x : std_logic_vector) return uint227_t is
  variable rv : uint227_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int227_t_to_slv(x : int227_t) return std_logic_vector is
  variable rv : std_logic_vector(226 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int227_t(x : std_logic_vector) return int227_t is
  variable rv : int227_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint228_t_to_slv(x : uint228_t) return std_logic_vector is
  variable rv : std_logic_vector(227 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint228_t(x : std_logic_vector) return uint228_t is
  variable rv : uint228_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int228_t_to_slv(x : int228_t) return std_logic_vector is
  variable rv : std_logic_vector(227 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int228_t(x : std_logic_vector) return int228_t is
  variable rv : int228_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint229_t_to_slv(x : uint229_t) return std_logic_vector is
  variable rv : std_logic_vector(228 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint229_t(x : std_logic_vector) return uint229_t is
  variable rv : uint229_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int229_t_to_slv(x : int229_t) return std_logic_vector is
  variable rv : std_logic_vector(228 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int229_t(x : std_logic_vector) return int229_t is
  variable rv : int229_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint230_t_to_slv(x : uint230_t) return std_logic_vector is
  variable rv : std_logic_vector(229 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint230_t(x : std_logic_vector) return uint230_t is
  variable rv : uint230_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int230_t_to_slv(x : int230_t) return std_logic_vector is
  variable rv : std_logic_vector(229 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int230_t(x : std_logic_vector) return int230_t is
  variable rv : int230_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint231_t_to_slv(x : uint231_t) return std_logic_vector is
  variable rv : std_logic_vector(230 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint231_t(x : std_logic_vector) return uint231_t is
  variable rv : uint231_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int231_t_to_slv(x : int231_t) return std_logic_vector is
  variable rv : std_logic_vector(230 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int231_t(x : std_logic_vector) return int231_t is
  variable rv : int231_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint232_t_to_slv(x : uint232_t) return std_logic_vector is
  variable rv : std_logic_vector(231 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint232_t(x : std_logic_vector) return uint232_t is
  variable rv : uint232_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int232_t_to_slv(x : int232_t) return std_logic_vector is
  variable rv : std_logic_vector(231 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int232_t(x : std_logic_vector) return int232_t is
  variable rv : int232_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint233_t_to_slv(x : uint233_t) return std_logic_vector is
  variable rv : std_logic_vector(232 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint233_t(x : std_logic_vector) return uint233_t is
  variable rv : uint233_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int233_t_to_slv(x : int233_t) return std_logic_vector is
  variable rv : std_logic_vector(232 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int233_t(x : std_logic_vector) return int233_t is
  variable rv : int233_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint234_t_to_slv(x : uint234_t) return std_logic_vector is
  variable rv : std_logic_vector(233 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint234_t(x : std_logic_vector) return uint234_t is
  variable rv : uint234_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int234_t_to_slv(x : int234_t) return std_logic_vector is
  variable rv : std_logic_vector(233 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int234_t(x : std_logic_vector) return int234_t is
  variable rv : int234_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint235_t_to_slv(x : uint235_t) return std_logic_vector is
  variable rv : std_logic_vector(234 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint235_t(x : std_logic_vector) return uint235_t is
  variable rv : uint235_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int235_t_to_slv(x : int235_t) return std_logic_vector is
  variable rv : std_logic_vector(234 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int235_t(x : std_logic_vector) return int235_t is
  variable rv : int235_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint236_t_to_slv(x : uint236_t) return std_logic_vector is
  variable rv : std_logic_vector(235 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint236_t(x : std_logic_vector) return uint236_t is
  variable rv : uint236_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int236_t_to_slv(x : int236_t) return std_logic_vector is
  variable rv : std_logic_vector(235 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int236_t(x : std_logic_vector) return int236_t is
  variable rv : int236_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint237_t_to_slv(x : uint237_t) return std_logic_vector is
  variable rv : std_logic_vector(236 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint237_t(x : std_logic_vector) return uint237_t is
  variable rv : uint237_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int237_t_to_slv(x : int237_t) return std_logic_vector is
  variable rv : std_logic_vector(236 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int237_t(x : std_logic_vector) return int237_t is
  variable rv : int237_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint238_t_to_slv(x : uint238_t) return std_logic_vector is
  variable rv : std_logic_vector(237 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint238_t(x : std_logic_vector) return uint238_t is
  variable rv : uint238_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int238_t_to_slv(x : int238_t) return std_logic_vector is
  variable rv : std_logic_vector(237 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int238_t(x : std_logic_vector) return int238_t is
  variable rv : int238_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint239_t_to_slv(x : uint239_t) return std_logic_vector is
  variable rv : std_logic_vector(238 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint239_t(x : std_logic_vector) return uint239_t is
  variable rv : uint239_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int239_t_to_slv(x : int239_t) return std_logic_vector is
  variable rv : std_logic_vector(238 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int239_t(x : std_logic_vector) return int239_t is
  variable rv : int239_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint240_t_to_slv(x : uint240_t) return std_logic_vector is
  variable rv : std_logic_vector(239 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint240_t(x : std_logic_vector) return uint240_t is
  variable rv : uint240_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int240_t_to_slv(x : int240_t) return std_logic_vector is
  variable rv : std_logic_vector(239 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int240_t(x : std_logic_vector) return int240_t is
  variable rv : int240_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint241_t_to_slv(x : uint241_t) return std_logic_vector is
  variable rv : std_logic_vector(240 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint241_t(x : std_logic_vector) return uint241_t is
  variable rv : uint241_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int241_t_to_slv(x : int241_t) return std_logic_vector is
  variable rv : std_logic_vector(240 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int241_t(x : std_logic_vector) return int241_t is
  variable rv : int241_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint242_t_to_slv(x : uint242_t) return std_logic_vector is
  variable rv : std_logic_vector(241 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint242_t(x : std_logic_vector) return uint242_t is
  variable rv : uint242_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int242_t_to_slv(x : int242_t) return std_logic_vector is
  variable rv : std_logic_vector(241 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int242_t(x : std_logic_vector) return int242_t is
  variable rv : int242_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint243_t_to_slv(x : uint243_t) return std_logic_vector is
  variable rv : std_logic_vector(242 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint243_t(x : std_logic_vector) return uint243_t is
  variable rv : uint243_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int243_t_to_slv(x : int243_t) return std_logic_vector is
  variable rv : std_logic_vector(242 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int243_t(x : std_logic_vector) return int243_t is
  variable rv : int243_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint244_t_to_slv(x : uint244_t) return std_logic_vector is
  variable rv : std_logic_vector(243 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint244_t(x : std_logic_vector) return uint244_t is
  variable rv : uint244_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int244_t_to_slv(x : int244_t) return std_logic_vector is
  variable rv : std_logic_vector(243 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int244_t(x : std_logic_vector) return int244_t is
  variable rv : int244_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint245_t_to_slv(x : uint245_t) return std_logic_vector is
  variable rv : std_logic_vector(244 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint245_t(x : std_logic_vector) return uint245_t is
  variable rv : uint245_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int245_t_to_slv(x : int245_t) return std_logic_vector is
  variable rv : std_logic_vector(244 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int245_t(x : std_logic_vector) return int245_t is
  variable rv : int245_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint246_t_to_slv(x : uint246_t) return std_logic_vector is
  variable rv : std_logic_vector(245 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint246_t(x : std_logic_vector) return uint246_t is
  variable rv : uint246_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int246_t_to_slv(x : int246_t) return std_logic_vector is
  variable rv : std_logic_vector(245 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int246_t(x : std_logic_vector) return int246_t is
  variable rv : int246_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint247_t_to_slv(x : uint247_t) return std_logic_vector is
  variable rv : std_logic_vector(246 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint247_t(x : std_logic_vector) return uint247_t is
  variable rv : uint247_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int247_t_to_slv(x : int247_t) return std_logic_vector is
  variable rv : std_logic_vector(246 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int247_t(x : std_logic_vector) return int247_t is
  variable rv : int247_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint248_t_to_slv(x : uint248_t) return std_logic_vector is
  variable rv : std_logic_vector(247 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint248_t(x : std_logic_vector) return uint248_t is
  variable rv : uint248_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int248_t_to_slv(x : int248_t) return std_logic_vector is
  variable rv : std_logic_vector(247 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int248_t(x : std_logic_vector) return int248_t is
  variable rv : int248_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint249_t_to_slv(x : uint249_t) return std_logic_vector is
  variable rv : std_logic_vector(248 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint249_t(x : std_logic_vector) return uint249_t is
  variable rv : uint249_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int249_t_to_slv(x : int249_t) return std_logic_vector is
  variable rv : std_logic_vector(248 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int249_t(x : std_logic_vector) return int249_t is
  variable rv : int249_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint250_t_to_slv(x : uint250_t) return std_logic_vector is
  variable rv : std_logic_vector(249 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint250_t(x : std_logic_vector) return uint250_t is
  variable rv : uint250_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int250_t_to_slv(x : int250_t) return std_logic_vector is
  variable rv : std_logic_vector(249 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int250_t(x : std_logic_vector) return int250_t is
  variable rv : int250_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint251_t_to_slv(x : uint251_t) return std_logic_vector is
  variable rv : std_logic_vector(250 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint251_t(x : std_logic_vector) return uint251_t is
  variable rv : uint251_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int251_t_to_slv(x : int251_t) return std_logic_vector is
  variable rv : std_logic_vector(250 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int251_t(x : std_logic_vector) return int251_t is
  variable rv : int251_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint252_t_to_slv(x : uint252_t) return std_logic_vector is
  variable rv : std_logic_vector(251 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint252_t(x : std_logic_vector) return uint252_t is
  variable rv : uint252_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int252_t_to_slv(x : int252_t) return std_logic_vector is
  variable rv : std_logic_vector(251 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int252_t(x : std_logic_vector) return int252_t is
  variable rv : int252_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint253_t_to_slv(x : uint253_t) return std_logic_vector is
  variable rv : std_logic_vector(252 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint253_t(x : std_logic_vector) return uint253_t is
  variable rv : uint253_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int253_t_to_slv(x : int253_t) return std_logic_vector is
  variable rv : std_logic_vector(252 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int253_t(x : std_logic_vector) return int253_t is
  variable rv : int253_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint254_t_to_slv(x : uint254_t) return std_logic_vector is
  variable rv : std_logic_vector(253 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint254_t(x : std_logic_vector) return uint254_t is
  variable rv : uint254_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int254_t_to_slv(x : int254_t) return std_logic_vector is
  variable rv : std_logic_vector(253 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int254_t(x : std_logic_vector) return int254_t is
  variable rv : int254_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint255_t_to_slv(x : uint255_t) return std_logic_vector is
  variable rv : std_logic_vector(254 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint255_t(x : std_logic_vector) return uint255_t is
  variable rv : uint255_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int255_t_to_slv(x : int255_t) return std_logic_vector is
  variable rv : std_logic_vector(254 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int255_t(x : std_logic_vector) return int255_t is
  variable rv : int255_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint256_t_to_slv(x : uint256_t) return std_logic_vector is
  variable rv : std_logic_vector(255 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint256_t(x : std_logic_vector) return uint256_t is
  variable rv : uint256_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int256_t_to_slv(x : int256_t) return std_logic_vector is
  variable rv : std_logic_vector(255 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int256_t(x : std_logic_vector) return int256_t is
  variable rv : int256_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint257_t_to_slv(x : uint257_t) return std_logic_vector is
  variable rv : std_logic_vector(256 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint257_t(x : std_logic_vector) return uint257_t is
  variable rv : uint257_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int257_t_to_slv(x : int257_t) return std_logic_vector is
  variable rv : std_logic_vector(256 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int257_t(x : std_logic_vector) return int257_t is
  variable rv : int257_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint258_t_to_slv(x : uint258_t) return std_logic_vector is
  variable rv : std_logic_vector(257 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint258_t(x : std_logic_vector) return uint258_t is
  variable rv : uint258_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int258_t_to_slv(x : int258_t) return std_logic_vector is
  variable rv : std_logic_vector(257 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int258_t(x : std_logic_vector) return int258_t is
  variable rv : int258_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint259_t_to_slv(x : uint259_t) return std_logic_vector is
  variable rv : std_logic_vector(258 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint259_t(x : std_logic_vector) return uint259_t is
  variable rv : uint259_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int259_t_to_slv(x : int259_t) return std_logic_vector is
  variable rv : std_logic_vector(258 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int259_t(x : std_logic_vector) return int259_t is
  variable rv : int259_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint260_t_to_slv(x : uint260_t) return std_logic_vector is
  variable rv : std_logic_vector(259 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint260_t(x : std_logic_vector) return uint260_t is
  variable rv : uint260_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int260_t_to_slv(x : int260_t) return std_logic_vector is
  variable rv : std_logic_vector(259 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int260_t(x : std_logic_vector) return int260_t is
  variable rv : int260_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint261_t_to_slv(x : uint261_t) return std_logic_vector is
  variable rv : std_logic_vector(260 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint261_t(x : std_logic_vector) return uint261_t is
  variable rv : uint261_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int261_t_to_slv(x : int261_t) return std_logic_vector is
  variable rv : std_logic_vector(260 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int261_t(x : std_logic_vector) return int261_t is
  variable rv : int261_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint262_t_to_slv(x : uint262_t) return std_logic_vector is
  variable rv : std_logic_vector(261 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint262_t(x : std_logic_vector) return uint262_t is
  variable rv : uint262_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int262_t_to_slv(x : int262_t) return std_logic_vector is
  variable rv : std_logic_vector(261 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int262_t(x : std_logic_vector) return int262_t is
  variable rv : int262_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint263_t_to_slv(x : uint263_t) return std_logic_vector is
  variable rv : std_logic_vector(262 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint263_t(x : std_logic_vector) return uint263_t is
  variable rv : uint263_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int263_t_to_slv(x : int263_t) return std_logic_vector is
  variable rv : std_logic_vector(262 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int263_t(x : std_logic_vector) return int263_t is
  variable rv : int263_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint264_t_to_slv(x : uint264_t) return std_logic_vector is
  variable rv : std_logic_vector(263 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint264_t(x : std_logic_vector) return uint264_t is
  variable rv : uint264_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int264_t_to_slv(x : int264_t) return std_logic_vector is
  variable rv : std_logic_vector(263 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int264_t(x : std_logic_vector) return int264_t is
  variable rv : int264_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint265_t_to_slv(x : uint265_t) return std_logic_vector is
  variable rv : std_logic_vector(264 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint265_t(x : std_logic_vector) return uint265_t is
  variable rv : uint265_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int265_t_to_slv(x : int265_t) return std_logic_vector is
  variable rv : std_logic_vector(264 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int265_t(x : std_logic_vector) return int265_t is
  variable rv : int265_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint266_t_to_slv(x : uint266_t) return std_logic_vector is
  variable rv : std_logic_vector(265 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint266_t(x : std_logic_vector) return uint266_t is
  variable rv : uint266_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int266_t_to_slv(x : int266_t) return std_logic_vector is
  variable rv : std_logic_vector(265 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int266_t(x : std_logic_vector) return int266_t is
  variable rv : int266_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint267_t_to_slv(x : uint267_t) return std_logic_vector is
  variable rv : std_logic_vector(266 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint267_t(x : std_logic_vector) return uint267_t is
  variable rv : uint267_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int267_t_to_slv(x : int267_t) return std_logic_vector is
  variable rv : std_logic_vector(266 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int267_t(x : std_logic_vector) return int267_t is
  variable rv : int267_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint268_t_to_slv(x : uint268_t) return std_logic_vector is
  variable rv : std_logic_vector(267 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint268_t(x : std_logic_vector) return uint268_t is
  variable rv : uint268_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int268_t_to_slv(x : int268_t) return std_logic_vector is
  variable rv : std_logic_vector(267 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int268_t(x : std_logic_vector) return int268_t is
  variable rv : int268_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint269_t_to_slv(x : uint269_t) return std_logic_vector is
  variable rv : std_logic_vector(268 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint269_t(x : std_logic_vector) return uint269_t is
  variable rv : uint269_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int269_t_to_slv(x : int269_t) return std_logic_vector is
  variable rv : std_logic_vector(268 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int269_t(x : std_logic_vector) return int269_t is
  variable rv : int269_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint270_t_to_slv(x : uint270_t) return std_logic_vector is
  variable rv : std_logic_vector(269 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint270_t(x : std_logic_vector) return uint270_t is
  variable rv : uint270_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int270_t_to_slv(x : int270_t) return std_logic_vector is
  variable rv : std_logic_vector(269 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int270_t(x : std_logic_vector) return int270_t is
  variable rv : int270_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint271_t_to_slv(x : uint271_t) return std_logic_vector is
  variable rv : std_logic_vector(270 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint271_t(x : std_logic_vector) return uint271_t is
  variable rv : uint271_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int271_t_to_slv(x : int271_t) return std_logic_vector is
  variable rv : std_logic_vector(270 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int271_t(x : std_logic_vector) return int271_t is
  variable rv : int271_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint272_t_to_slv(x : uint272_t) return std_logic_vector is
  variable rv : std_logic_vector(271 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint272_t(x : std_logic_vector) return uint272_t is
  variable rv : uint272_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int272_t_to_slv(x : int272_t) return std_logic_vector is
  variable rv : std_logic_vector(271 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int272_t(x : std_logic_vector) return int272_t is
  variable rv : int272_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint273_t_to_slv(x : uint273_t) return std_logic_vector is
  variable rv : std_logic_vector(272 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint273_t(x : std_logic_vector) return uint273_t is
  variable rv : uint273_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int273_t_to_slv(x : int273_t) return std_logic_vector is
  variable rv : std_logic_vector(272 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int273_t(x : std_logic_vector) return int273_t is
  variable rv : int273_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint274_t_to_slv(x : uint274_t) return std_logic_vector is
  variable rv : std_logic_vector(273 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint274_t(x : std_logic_vector) return uint274_t is
  variable rv : uint274_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int274_t_to_slv(x : int274_t) return std_logic_vector is
  variable rv : std_logic_vector(273 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int274_t(x : std_logic_vector) return int274_t is
  variable rv : int274_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint275_t_to_slv(x : uint275_t) return std_logic_vector is
  variable rv : std_logic_vector(274 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint275_t(x : std_logic_vector) return uint275_t is
  variable rv : uint275_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int275_t_to_slv(x : int275_t) return std_logic_vector is
  variable rv : std_logic_vector(274 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int275_t(x : std_logic_vector) return int275_t is
  variable rv : int275_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint276_t_to_slv(x : uint276_t) return std_logic_vector is
  variable rv : std_logic_vector(275 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint276_t(x : std_logic_vector) return uint276_t is
  variable rv : uint276_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int276_t_to_slv(x : int276_t) return std_logic_vector is
  variable rv : std_logic_vector(275 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int276_t(x : std_logic_vector) return int276_t is
  variable rv : int276_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint277_t_to_slv(x : uint277_t) return std_logic_vector is
  variable rv : std_logic_vector(276 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint277_t(x : std_logic_vector) return uint277_t is
  variable rv : uint277_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int277_t_to_slv(x : int277_t) return std_logic_vector is
  variable rv : std_logic_vector(276 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int277_t(x : std_logic_vector) return int277_t is
  variable rv : int277_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint278_t_to_slv(x : uint278_t) return std_logic_vector is
  variable rv : std_logic_vector(277 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint278_t(x : std_logic_vector) return uint278_t is
  variable rv : uint278_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int278_t_to_slv(x : int278_t) return std_logic_vector is
  variable rv : std_logic_vector(277 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int278_t(x : std_logic_vector) return int278_t is
  variable rv : int278_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint279_t_to_slv(x : uint279_t) return std_logic_vector is
  variable rv : std_logic_vector(278 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint279_t(x : std_logic_vector) return uint279_t is
  variable rv : uint279_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int279_t_to_slv(x : int279_t) return std_logic_vector is
  variable rv : std_logic_vector(278 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int279_t(x : std_logic_vector) return int279_t is
  variable rv : int279_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint280_t_to_slv(x : uint280_t) return std_logic_vector is
  variable rv : std_logic_vector(279 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint280_t(x : std_logic_vector) return uint280_t is
  variable rv : uint280_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int280_t_to_slv(x : int280_t) return std_logic_vector is
  variable rv : std_logic_vector(279 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int280_t(x : std_logic_vector) return int280_t is
  variable rv : int280_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint281_t_to_slv(x : uint281_t) return std_logic_vector is
  variable rv : std_logic_vector(280 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint281_t(x : std_logic_vector) return uint281_t is
  variable rv : uint281_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int281_t_to_slv(x : int281_t) return std_logic_vector is
  variable rv : std_logic_vector(280 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int281_t(x : std_logic_vector) return int281_t is
  variable rv : int281_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint282_t_to_slv(x : uint282_t) return std_logic_vector is
  variable rv : std_logic_vector(281 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint282_t(x : std_logic_vector) return uint282_t is
  variable rv : uint282_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int282_t_to_slv(x : int282_t) return std_logic_vector is
  variable rv : std_logic_vector(281 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int282_t(x : std_logic_vector) return int282_t is
  variable rv : int282_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint283_t_to_slv(x : uint283_t) return std_logic_vector is
  variable rv : std_logic_vector(282 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint283_t(x : std_logic_vector) return uint283_t is
  variable rv : uint283_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int283_t_to_slv(x : int283_t) return std_logic_vector is
  variable rv : std_logic_vector(282 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int283_t(x : std_logic_vector) return int283_t is
  variable rv : int283_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint284_t_to_slv(x : uint284_t) return std_logic_vector is
  variable rv : std_logic_vector(283 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint284_t(x : std_logic_vector) return uint284_t is
  variable rv : uint284_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int284_t_to_slv(x : int284_t) return std_logic_vector is
  variable rv : std_logic_vector(283 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int284_t(x : std_logic_vector) return int284_t is
  variable rv : int284_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint285_t_to_slv(x : uint285_t) return std_logic_vector is
  variable rv : std_logic_vector(284 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint285_t(x : std_logic_vector) return uint285_t is
  variable rv : uint285_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int285_t_to_slv(x : int285_t) return std_logic_vector is
  variable rv : std_logic_vector(284 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int285_t(x : std_logic_vector) return int285_t is
  variable rv : int285_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint286_t_to_slv(x : uint286_t) return std_logic_vector is
  variable rv : std_logic_vector(285 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint286_t(x : std_logic_vector) return uint286_t is
  variable rv : uint286_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int286_t_to_slv(x : int286_t) return std_logic_vector is
  variable rv : std_logic_vector(285 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int286_t(x : std_logic_vector) return int286_t is
  variable rv : int286_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint287_t_to_slv(x : uint287_t) return std_logic_vector is
  variable rv : std_logic_vector(286 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint287_t(x : std_logic_vector) return uint287_t is
  variable rv : uint287_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int287_t_to_slv(x : int287_t) return std_logic_vector is
  variable rv : std_logic_vector(286 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int287_t(x : std_logic_vector) return int287_t is
  variable rv : int287_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint288_t_to_slv(x : uint288_t) return std_logic_vector is
  variable rv : std_logic_vector(287 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint288_t(x : std_logic_vector) return uint288_t is
  variable rv : uint288_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int288_t_to_slv(x : int288_t) return std_logic_vector is
  variable rv : std_logic_vector(287 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int288_t(x : std_logic_vector) return int288_t is
  variable rv : int288_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint289_t_to_slv(x : uint289_t) return std_logic_vector is
  variable rv : std_logic_vector(288 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint289_t(x : std_logic_vector) return uint289_t is
  variable rv : uint289_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int289_t_to_slv(x : int289_t) return std_logic_vector is
  variable rv : std_logic_vector(288 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int289_t(x : std_logic_vector) return int289_t is
  variable rv : int289_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint290_t_to_slv(x : uint290_t) return std_logic_vector is
  variable rv : std_logic_vector(289 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint290_t(x : std_logic_vector) return uint290_t is
  variable rv : uint290_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int290_t_to_slv(x : int290_t) return std_logic_vector is
  variable rv : std_logic_vector(289 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int290_t(x : std_logic_vector) return int290_t is
  variable rv : int290_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint291_t_to_slv(x : uint291_t) return std_logic_vector is
  variable rv : std_logic_vector(290 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint291_t(x : std_logic_vector) return uint291_t is
  variable rv : uint291_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int291_t_to_slv(x : int291_t) return std_logic_vector is
  variable rv : std_logic_vector(290 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int291_t(x : std_logic_vector) return int291_t is
  variable rv : int291_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint292_t_to_slv(x : uint292_t) return std_logic_vector is
  variable rv : std_logic_vector(291 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint292_t(x : std_logic_vector) return uint292_t is
  variable rv : uint292_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int292_t_to_slv(x : int292_t) return std_logic_vector is
  variable rv : std_logic_vector(291 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int292_t(x : std_logic_vector) return int292_t is
  variable rv : int292_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint293_t_to_slv(x : uint293_t) return std_logic_vector is
  variable rv : std_logic_vector(292 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint293_t(x : std_logic_vector) return uint293_t is
  variable rv : uint293_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int293_t_to_slv(x : int293_t) return std_logic_vector is
  variable rv : std_logic_vector(292 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int293_t(x : std_logic_vector) return int293_t is
  variable rv : int293_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint294_t_to_slv(x : uint294_t) return std_logic_vector is
  variable rv : std_logic_vector(293 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint294_t(x : std_logic_vector) return uint294_t is
  variable rv : uint294_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int294_t_to_slv(x : int294_t) return std_logic_vector is
  variable rv : std_logic_vector(293 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int294_t(x : std_logic_vector) return int294_t is
  variable rv : int294_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint295_t_to_slv(x : uint295_t) return std_logic_vector is
  variable rv : std_logic_vector(294 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint295_t(x : std_logic_vector) return uint295_t is
  variable rv : uint295_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int295_t_to_slv(x : int295_t) return std_logic_vector is
  variable rv : std_logic_vector(294 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int295_t(x : std_logic_vector) return int295_t is
  variable rv : int295_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint296_t_to_slv(x : uint296_t) return std_logic_vector is
  variable rv : std_logic_vector(295 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint296_t(x : std_logic_vector) return uint296_t is
  variable rv : uint296_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int296_t_to_slv(x : int296_t) return std_logic_vector is
  variable rv : std_logic_vector(295 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int296_t(x : std_logic_vector) return int296_t is
  variable rv : int296_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint297_t_to_slv(x : uint297_t) return std_logic_vector is
  variable rv : std_logic_vector(296 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint297_t(x : std_logic_vector) return uint297_t is
  variable rv : uint297_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int297_t_to_slv(x : int297_t) return std_logic_vector is
  variable rv : std_logic_vector(296 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int297_t(x : std_logic_vector) return int297_t is
  variable rv : int297_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint298_t_to_slv(x : uint298_t) return std_logic_vector is
  variable rv : std_logic_vector(297 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint298_t(x : std_logic_vector) return uint298_t is
  variable rv : uint298_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int298_t_to_slv(x : int298_t) return std_logic_vector is
  variable rv : std_logic_vector(297 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int298_t(x : std_logic_vector) return int298_t is
  variable rv : int298_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint299_t_to_slv(x : uint299_t) return std_logic_vector is
  variable rv : std_logic_vector(298 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint299_t(x : std_logic_vector) return uint299_t is
  variable rv : uint299_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int299_t_to_slv(x : int299_t) return std_logic_vector is
  variable rv : std_logic_vector(298 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int299_t(x : std_logic_vector) return int299_t is
  variable rv : int299_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint300_t_to_slv(x : uint300_t) return std_logic_vector is
  variable rv : std_logic_vector(299 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint300_t(x : std_logic_vector) return uint300_t is
  variable rv : uint300_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int300_t_to_slv(x : int300_t) return std_logic_vector is
  variable rv : std_logic_vector(299 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int300_t(x : std_logic_vector) return int300_t is
  variable rv : int300_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint301_t_to_slv(x : uint301_t) return std_logic_vector is
  variable rv : std_logic_vector(300 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint301_t(x : std_logic_vector) return uint301_t is
  variable rv : uint301_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int301_t_to_slv(x : int301_t) return std_logic_vector is
  variable rv : std_logic_vector(300 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int301_t(x : std_logic_vector) return int301_t is
  variable rv : int301_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint302_t_to_slv(x : uint302_t) return std_logic_vector is
  variable rv : std_logic_vector(301 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint302_t(x : std_logic_vector) return uint302_t is
  variable rv : uint302_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int302_t_to_slv(x : int302_t) return std_logic_vector is
  variable rv : std_logic_vector(301 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int302_t(x : std_logic_vector) return int302_t is
  variable rv : int302_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint303_t_to_slv(x : uint303_t) return std_logic_vector is
  variable rv : std_logic_vector(302 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint303_t(x : std_logic_vector) return uint303_t is
  variable rv : uint303_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int303_t_to_slv(x : int303_t) return std_logic_vector is
  variable rv : std_logic_vector(302 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int303_t(x : std_logic_vector) return int303_t is
  variable rv : int303_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint304_t_to_slv(x : uint304_t) return std_logic_vector is
  variable rv : std_logic_vector(303 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint304_t(x : std_logic_vector) return uint304_t is
  variable rv : uint304_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int304_t_to_slv(x : int304_t) return std_logic_vector is
  variable rv : std_logic_vector(303 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int304_t(x : std_logic_vector) return int304_t is
  variable rv : int304_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint305_t_to_slv(x : uint305_t) return std_logic_vector is
  variable rv : std_logic_vector(304 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint305_t(x : std_logic_vector) return uint305_t is
  variable rv : uint305_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int305_t_to_slv(x : int305_t) return std_logic_vector is
  variable rv : std_logic_vector(304 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int305_t(x : std_logic_vector) return int305_t is
  variable rv : int305_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint306_t_to_slv(x : uint306_t) return std_logic_vector is
  variable rv : std_logic_vector(305 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint306_t(x : std_logic_vector) return uint306_t is
  variable rv : uint306_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int306_t_to_slv(x : int306_t) return std_logic_vector is
  variable rv : std_logic_vector(305 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int306_t(x : std_logic_vector) return int306_t is
  variable rv : int306_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint307_t_to_slv(x : uint307_t) return std_logic_vector is
  variable rv : std_logic_vector(306 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint307_t(x : std_logic_vector) return uint307_t is
  variable rv : uint307_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int307_t_to_slv(x : int307_t) return std_logic_vector is
  variable rv : std_logic_vector(306 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int307_t(x : std_logic_vector) return int307_t is
  variable rv : int307_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint308_t_to_slv(x : uint308_t) return std_logic_vector is
  variable rv : std_logic_vector(307 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint308_t(x : std_logic_vector) return uint308_t is
  variable rv : uint308_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int308_t_to_slv(x : int308_t) return std_logic_vector is
  variable rv : std_logic_vector(307 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int308_t(x : std_logic_vector) return int308_t is
  variable rv : int308_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint309_t_to_slv(x : uint309_t) return std_logic_vector is
  variable rv : std_logic_vector(308 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint309_t(x : std_logic_vector) return uint309_t is
  variable rv : uint309_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int309_t_to_slv(x : int309_t) return std_logic_vector is
  variable rv : std_logic_vector(308 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int309_t(x : std_logic_vector) return int309_t is
  variable rv : int309_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint310_t_to_slv(x : uint310_t) return std_logic_vector is
  variable rv : std_logic_vector(309 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint310_t(x : std_logic_vector) return uint310_t is
  variable rv : uint310_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int310_t_to_slv(x : int310_t) return std_logic_vector is
  variable rv : std_logic_vector(309 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int310_t(x : std_logic_vector) return int310_t is
  variable rv : int310_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint311_t_to_slv(x : uint311_t) return std_logic_vector is
  variable rv : std_logic_vector(310 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint311_t(x : std_logic_vector) return uint311_t is
  variable rv : uint311_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int311_t_to_slv(x : int311_t) return std_logic_vector is
  variable rv : std_logic_vector(310 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int311_t(x : std_logic_vector) return int311_t is
  variable rv : int311_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint312_t_to_slv(x : uint312_t) return std_logic_vector is
  variable rv : std_logic_vector(311 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint312_t(x : std_logic_vector) return uint312_t is
  variable rv : uint312_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int312_t_to_slv(x : int312_t) return std_logic_vector is
  variable rv : std_logic_vector(311 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int312_t(x : std_logic_vector) return int312_t is
  variable rv : int312_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint313_t_to_slv(x : uint313_t) return std_logic_vector is
  variable rv : std_logic_vector(312 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint313_t(x : std_logic_vector) return uint313_t is
  variable rv : uint313_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int313_t_to_slv(x : int313_t) return std_logic_vector is
  variable rv : std_logic_vector(312 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int313_t(x : std_logic_vector) return int313_t is
  variable rv : int313_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint314_t_to_slv(x : uint314_t) return std_logic_vector is
  variable rv : std_logic_vector(313 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint314_t(x : std_logic_vector) return uint314_t is
  variable rv : uint314_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int314_t_to_slv(x : int314_t) return std_logic_vector is
  variable rv : std_logic_vector(313 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int314_t(x : std_logic_vector) return int314_t is
  variable rv : int314_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint315_t_to_slv(x : uint315_t) return std_logic_vector is
  variable rv : std_logic_vector(314 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint315_t(x : std_logic_vector) return uint315_t is
  variable rv : uint315_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int315_t_to_slv(x : int315_t) return std_logic_vector is
  variable rv : std_logic_vector(314 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int315_t(x : std_logic_vector) return int315_t is
  variable rv : int315_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint316_t_to_slv(x : uint316_t) return std_logic_vector is
  variable rv : std_logic_vector(315 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint316_t(x : std_logic_vector) return uint316_t is
  variable rv : uint316_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int316_t_to_slv(x : int316_t) return std_logic_vector is
  variable rv : std_logic_vector(315 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int316_t(x : std_logic_vector) return int316_t is
  variable rv : int316_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint317_t_to_slv(x : uint317_t) return std_logic_vector is
  variable rv : std_logic_vector(316 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint317_t(x : std_logic_vector) return uint317_t is
  variable rv : uint317_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int317_t_to_slv(x : int317_t) return std_logic_vector is
  variable rv : std_logic_vector(316 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int317_t(x : std_logic_vector) return int317_t is
  variable rv : int317_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint318_t_to_slv(x : uint318_t) return std_logic_vector is
  variable rv : std_logic_vector(317 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint318_t(x : std_logic_vector) return uint318_t is
  variable rv : uint318_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int318_t_to_slv(x : int318_t) return std_logic_vector is
  variable rv : std_logic_vector(317 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int318_t(x : std_logic_vector) return int318_t is
  variable rv : int318_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint319_t_to_slv(x : uint319_t) return std_logic_vector is
  variable rv : std_logic_vector(318 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint319_t(x : std_logic_vector) return uint319_t is
  variable rv : uint319_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int319_t_to_slv(x : int319_t) return std_logic_vector is
  variable rv : std_logic_vector(318 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int319_t(x : std_logic_vector) return int319_t is
  variable rv : int319_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint320_t_to_slv(x : uint320_t) return std_logic_vector is
  variable rv : std_logic_vector(319 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint320_t(x : std_logic_vector) return uint320_t is
  variable rv : uint320_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int320_t_to_slv(x : int320_t) return std_logic_vector is
  variable rv : std_logic_vector(319 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int320_t(x : std_logic_vector) return int320_t is
  variable rv : int320_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint321_t_to_slv(x : uint321_t) return std_logic_vector is
  variable rv : std_logic_vector(320 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint321_t(x : std_logic_vector) return uint321_t is
  variable rv : uint321_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int321_t_to_slv(x : int321_t) return std_logic_vector is
  variable rv : std_logic_vector(320 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int321_t(x : std_logic_vector) return int321_t is
  variable rv : int321_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint322_t_to_slv(x : uint322_t) return std_logic_vector is
  variable rv : std_logic_vector(321 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint322_t(x : std_logic_vector) return uint322_t is
  variable rv : uint322_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int322_t_to_slv(x : int322_t) return std_logic_vector is
  variable rv : std_logic_vector(321 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int322_t(x : std_logic_vector) return int322_t is
  variable rv : int322_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint323_t_to_slv(x : uint323_t) return std_logic_vector is
  variable rv : std_logic_vector(322 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint323_t(x : std_logic_vector) return uint323_t is
  variable rv : uint323_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int323_t_to_slv(x : int323_t) return std_logic_vector is
  variable rv : std_logic_vector(322 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int323_t(x : std_logic_vector) return int323_t is
  variable rv : int323_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint324_t_to_slv(x : uint324_t) return std_logic_vector is
  variable rv : std_logic_vector(323 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint324_t(x : std_logic_vector) return uint324_t is
  variable rv : uint324_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int324_t_to_slv(x : int324_t) return std_logic_vector is
  variable rv : std_logic_vector(323 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int324_t(x : std_logic_vector) return int324_t is
  variable rv : int324_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint325_t_to_slv(x : uint325_t) return std_logic_vector is
  variable rv : std_logic_vector(324 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint325_t(x : std_logic_vector) return uint325_t is
  variable rv : uint325_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int325_t_to_slv(x : int325_t) return std_logic_vector is
  variable rv : std_logic_vector(324 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int325_t(x : std_logic_vector) return int325_t is
  variable rv : int325_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint326_t_to_slv(x : uint326_t) return std_logic_vector is
  variable rv : std_logic_vector(325 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint326_t(x : std_logic_vector) return uint326_t is
  variable rv : uint326_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int326_t_to_slv(x : int326_t) return std_logic_vector is
  variable rv : std_logic_vector(325 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int326_t(x : std_logic_vector) return int326_t is
  variable rv : int326_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint327_t_to_slv(x : uint327_t) return std_logic_vector is
  variable rv : std_logic_vector(326 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint327_t(x : std_logic_vector) return uint327_t is
  variable rv : uint327_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int327_t_to_slv(x : int327_t) return std_logic_vector is
  variable rv : std_logic_vector(326 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int327_t(x : std_logic_vector) return int327_t is
  variable rv : int327_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint328_t_to_slv(x : uint328_t) return std_logic_vector is
  variable rv : std_logic_vector(327 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint328_t(x : std_logic_vector) return uint328_t is
  variable rv : uint328_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int328_t_to_slv(x : int328_t) return std_logic_vector is
  variable rv : std_logic_vector(327 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int328_t(x : std_logic_vector) return int328_t is
  variable rv : int328_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint329_t_to_slv(x : uint329_t) return std_logic_vector is
  variable rv : std_logic_vector(328 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint329_t(x : std_logic_vector) return uint329_t is
  variable rv : uint329_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int329_t_to_slv(x : int329_t) return std_logic_vector is
  variable rv : std_logic_vector(328 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int329_t(x : std_logic_vector) return int329_t is
  variable rv : int329_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint330_t_to_slv(x : uint330_t) return std_logic_vector is
  variable rv : std_logic_vector(329 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint330_t(x : std_logic_vector) return uint330_t is
  variable rv : uint330_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int330_t_to_slv(x : int330_t) return std_logic_vector is
  variable rv : std_logic_vector(329 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int330_t(x : std_logic_vector) return int330_t is
  variable rv : int330_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint331_t_to_slv(x : uint331_t) return std_logic_vector is
  variable rv : std_logic_vector(330 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint331_t(x : std_logic_vector) return uint331_t is
  variable rv : uint331_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int331_t_to_slv(x : int331_t) return std_logic_vector is
  variable rv : std_logic_vector(330 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int331_t(x : std_logic_vector) return int331_t is
  variable rv : int331_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint332_t_to_slv(x : uint332_t) return std_logic_vector is
  variable rv : std_logic_vector(331 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint332_t(x : std_logic_vector) return uint332_t is
  variable rv : uint332_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int332_t_to_slv(x : int332_t) return std_logic_vector is
  variable rv : std_logic_vector(331 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int332_t(x : std_logic_vector) return int332_t is
  variable rv : int332_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint333_t_to_slv(x : uint333_t) return std_logic_vector is
  variable rv : std_logic_vector(332 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint333_t(x : std_logic_vector) return uint333_t is
  variable rv : uint333_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int333_t_to_slv(x : int333_t) return std_logic_vector is
  variable rv : std_logic_vector(332 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int333_t(x : std_logic_vector) return int333_t is
  variable rv : int333_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint334_t_to_slv(x : uint334_t) return std_logic_vector is
  variable rv : std_logic_vector(333 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint334_t(x : std_logic_vector) return uint334_t is
  variable rv : uint334_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int334_t_to_slv(x : int334_t) return std_logic_vector is
  variable rv : std_logic_vector(333 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int334_t(x : std_logic_vector) return int334_t is
  variable rv : int334_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint335_t_to_slv(x : uint335_t) return std_logic_vector is
  variable rv : std_logic_vector(334 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint335_t(x : std_logic_vector) return uint335_t is
  variable rv : uint335_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int335_t_to_slv(x : int335_t) return std_logic_vector is
  variable rv : std_logic_vector(334 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int335_t(x : std_logic_vector) return int335_t is
  variable rv : int335_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint336_t_to_slv(x : uint336_t) return std_logic_vector is
  variable rv : std_logic_vector(335 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint336_t(x : std_logic_vector) return uint336_t is
  variable rv : uint336_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int336_t_to_slv(x : int336_t) return std_logic_vector is
  variable rv : std_logic_vector(335 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int336_t(x : std_logic_vector) return int336_t is
  variable rv : int336_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint337_t_to_slv(x : uint337_t) return std_logic_vector is
  variable rv : std_logic_vector(336 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint337_t(x : std_logic_vector) return uint337_t is
  variable rv : uint337_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int337_t_to_slv(x : int337_t) return std_logic_vector is
  variable rv : std_logic_vector(336 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int337_t(x : std_logic_vector) return int337_t is
  variable rv : int337_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint338_t_to_slv(x : uint338_t) return std_logic_vector is
  variable rv : std_logic_vector(337 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint338_t(x : std_logic_vector) return uint338_t is
  variable rv : uint338_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int338_t_to_slv(x : int338_t) return std_logic_vector is
  variable rv : std_logic_vector(337 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int338_t(x : std_logic_vector) return int338_t is
  variable rv : int338_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint339_t_to_slv(x : uint339_t) return std_logic_vector is
  variable rv : std_logic_vector(338 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint339_t(x : std_logic_vector) return uint339_t is
  variable rv : uint339_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int339_t_to_slv(x : int339_t) return std_logic_vector is
  variable rv : std_logic_vector(338 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int339_t(x : std_logic_vector) return int339_t is
  variable rv : int339_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint340_t_to_slv(x : uint340_t) return std_logic_vector is
  variable rv : std_logic_vector(339 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint340_t(x : std_logic_vector) return uint340_t is
  variable rv : uint340_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int340_t_to_slv(x : int340_t) return std_logic_vector is
  variable rv : std_logic_vector(339 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int340_t(x : std_logic_vector) return int340_t is
  variable rv : int340_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint341_t_to_slv(x : uint341_t) return std_logic_vector is
  variable rv : std_logic_vector(340 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint341_t(x : std_logic_vector) return uint341_t is
  variable rv : uint341_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int341_t_to_slv(x : int341_t) return std_logic_vector is
  variable rv : std_logic_vector(340 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int341_t(x : std_logic_vector) return int341_t is
  variable rv : int341_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint342_t_to_slv(x : uint342_t) return std_logic_vector is
  variable rv : std_logic_vector(341 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint342_t(x : std_logic_vector) return uint342_t is
  variable rv : uint342_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int342_t_to_slv(x : int342_t) return std_logic_vector is
  variable rv : std_logic_vector(341 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int342_t(x : std_logic_vector) return int342_t is
  variable rv : int342_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint343_t_to_slv(x : uint343_t) return std_logic_vector is
  variable rv : std_logic_vector(342 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint343_t(x : std_logic_vector) return uint343_t is
  variable rv : uint343_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int343_t_to_slv(x : int343_t) return std_logic_vector is
  variable rv : std_logic_vector(342 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int343_t(x : std_logic_vector) return int343_t is
  variable rv : int343_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint344_t_to_slv(x : uint344_t) return std_logic_vector is
  variable rv : std_logic_vector(343 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint344_t(x : std_logic_vector) return uint344_t is
  variable rv : uint344_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int344_t_to_slv(x : int344_t) return std_logic_vector is
  variable rv : std_logic_vector(343 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int344_t(x : std_logic_vector) return int344_t is
  variable rv : int344_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint345_t_to_slv(x : uint345_t) return std_logic_vector is
  variable rv : std_logic_vector(344 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint345_t(x : std_logic_vector) return uint345_t is
  variable rv : uint345_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int345_t_to_slv(x : int345_t) return std_logic_vector is
  variable rv : std_logic_vector(344 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int345_t(x : std_logic_vector) return int345_t is
  variable rv : int345_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint346_t_to_slv(x : uint346_t) return std_logic_vector is
  variable rv : std_logic_vector(345 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint346_t(x : std_logic_vector) return uint346_t is
  variable rv : uint346_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int346_t_to_slv(x : int346_t) return std_logic_vector is
  variable rv : std_logic_vector(345 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int346_t(x : std_logic_vector) return int346_t is
  variable rv : int346_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint347_t_to_slv(x : uint347_t) return std_logic_vector is
  variable rv : std_logic_vector(346 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint347_t(x : std_logic_vector) return uint347_t is
  variable rv : uint347_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int347_t_to_slv(x : int347_t) return std_logic_vector is
  variable rv : std_logic_vector(346 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int347_t(x : std_logic_vector) return int347_t is
  variable rv : int347_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint348_t_to_slv(x : uint348_t) return std_logic_vector is
  variable rv : std_logic_vector(347 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint348_t(x : std_logic_vector) return uint348_t is
  variable rv : uint348_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int348_t_to_slv(x : int348_t) return std_logic_vector is
  variable rv : std_logic_vector(347 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int348_t(x : std_logic_vector) return int348_t is
  variable rv : int348_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint349_t_to_slv(x : uint349_t) return std_logic_vector is
  variable rv : std_logic_vector(348 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint349_t(x : std_logic_vector) return uint349_t is
  variable rv : uint349_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int349_t_to_slv(x : int349_t) return std_logic_vector is
  variable rv : std_logic_vector(348 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int349_t(x : std_logic_vector) return int349_t is
  variable rv : int349_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint350_t_to_slv(x : uint350_t) return std_logic_vector is
  variable rv : std_logic_vector(349 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint350_t(x : std_logic_vector) return uint350_t is
  variable rv : uint350_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int350_t_to_slv(x : int350_t) return std_logic_vector is
  variable rv : std_logic_vector(349 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int350_t(x : std_logic_vector) return int350_t is
  variable rv : int350_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint351_t_to_slv(x : uint351_t) return std_logic_vector is
  variable rv : std_logic_vector(350 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint351_t(x : std_logic_vector) return uint351_t is
  variable rv : uint351_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int351_t_to_slv(x : int351_t) return std_logic_vector is
  variable rv : std_logic_vector(350 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int351_t(x : std_logic_vector) return int351_t is
  variable rv : int351_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint352_t_to_slv(x : uint352_t) return std_logic_vector is
  variable rv : std_logic_vector(351 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint352_t(x : std_logic_vector) return uint352_t is
  variable rv : uint352_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int352_t_to_slv(x : int352_t) return std_logic_vector is
  variable rv : std_logic_vector(351 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int352_t(x : std_logic_vector) return int352_t is
  variable rv : int352_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint353_t_to_slv(x : uint353_t) return std_logic_vector is
  variable rv : std_logic_vector(352 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint353_t(x : std_logic_vector) return uint353_t is
  variable rv : uint353_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int353_t_to_slv(x : int353_t) return std_logic_vector is
  variable rv : std_logic_vector(352 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int353_t(x : std_logic_vector) return int353_t is
  variable rv : int353_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint354_t_to_slv(x : uint354_t) return std_logic_vector is
  variable rv : std_logic_vector(353 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint354_t(x : std_logic_vector) return uint354_t is
  variable rv : uint354_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int354_t_to_slv(x : int354_t) return std_logic_vector is
  variable rv : std_logic_vector(353 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int354_t(x : std_logic_vector) return int354_t is
  variable rv : int354_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint355_t_to_slv(x : uint355_t) return std_logic_vector is
  variable rv : std_logic_vector(354 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint355_t(x : std_logic_vector) return uint355_t is
  variable rv : uint355_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int355_t_to_slv(x : int355_t) return std_logic_vector is
  variable rv : std_logic_vector(354 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int355_t(x : std_logic_vector) return int355_t is
  variable rv : int355_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint356_t_to_slv(x : uint356_t) return std_logic_vector is
  variable rv : std_logic_vector(355 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint356_t(x : std_logic_vector) return uint356_t is
  variable rv : uint356_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int356_t_to_slv(x : int356_t) return std_logic_vector is
  variable rv : std_logic_vector(355 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int356_t(x : std_logic_vector) return int356_t is
  variable rv : int356_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint357_t_to_slv(x : uint357_t) return std_logic_vector is
  variable rv : std_logic_vector(356 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint357_t(x : std_logic_vector) return uint357_t is
  variable rv : uint357_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int357_t_to_slv(x : int357_t) return std_logic_vector is
  variable rv : std_logic_vector(356 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int357_t(x : std_logic_vector) return int357_t is
  variable rv : int357_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint358_t_to_slv(x : uint358_t) return std_logic_vector is
  variable rv : std_logic_vector(357 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint358_t(x : std_logic_vector) return uint358_t is
  variable rv : uint358_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int358_t_to_slv(x : int358_t) return std_logic_vector is
  variable rv : std_logic_vector(357 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int358_t(x : std_logic_vector) return int358_t is
  variable rv : int358_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint359_t_to_slv(x : uint359_t) return std_logic_vector is
  variable rv : std_logic_vector(358 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint359_t(x : std_logic_vector) return uint359_t is
  variable rv : uint359_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int359_t_to_slv(x : int359_t) return std_logic_vector is
  variable rv : std_logic_vector(358 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int359_t(x : std_logic_vector) return int359_t is
  variable rv : int359_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint360_t_to_slv(x : uint360_t) return std_logic_vector is
  variable rv : std_logic_vector(359 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint360_t(x : std_logic_vector) return uint360_t is
  variable rv : uint360_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int360_t_to_slv(x : int360_t) return std_logic_vector is
  variable rv : std_logic_vector(359 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int360_t(x : std_logic_vector) return int360_t is
  variable rv : int360_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint361_t_to_slv(x : uint361_t) return std_logic_vector is
  variable rv : std_logic_vector(360 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint361_t(x : std_logic_vector) return uint361_t is
  variable rv : uint361_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int361_t_to_slv(x : int361_t) return std_logic_vector is
  variable rv : std_logic_vector(360 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int361_t(x : std_logic_vector) return int361_t is
  variable rv : int361_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint362_t_to_slv(x : uint362_t) return std_logic_vector is
  variable rv : std_logic_vector(361 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint362_t(x : std_logic_vector) return uint362_t is
  variable rv : uint362_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int362_t_to_slv(x : int362_t) return std_logic_vector is
  variable rv : std_logic_vector(361 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int362_t(x : std_logic_vector) return int362_t is
  variable rv : int362_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint363_t_to_slv(x : uint363_t) return std_logic_vector is
  variable rv : std_logic_vector(362 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint363_t(x : std_logic_vector) return uint363_t is
  variable rv : uint363_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int363_t_to_slv(x : int363_t) return std_logic_vector is
  variable rv : std_logic_vector(362 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int363_t(x : std_logic_vector) return int363_t is
  variable rv : int363_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint364_t_to_slv(x : uint364_t) return std_logic_vector is
  variable rv : std_logic_vector(363 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint364_t(x : std_logic_vector) return uint364_t is
  variable rv : uint364_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int364_t_to_slv(x : int364_t) return std_logic_vector is
  variable rv : std_logic_vector(363 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int364_t(x : std_logic_vector) return int364_t is
  variable rv : int364_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint365_t_to_slv(x : uint365_t) return std_logic_vector is
  variable rv : std_logic_vector(364 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint365_t(x : std_logic_vector) return uint365_t is
  variable rv : uint365_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int365_t_to_slv(x : int365_t) return std_logic_vector is
  variable rv : std_logic_vector(364 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int365_t(x : std_logic_vector) return int365_t is
  variable rv : int365_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint366_t_to_slv(x : uint366_t) return std_logic_vector is
  variable rv : std_logic_vector(365 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint366_t(x : std_logic_vector) return uint366_t is
  variable rv : uint366_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int366_t_to_slv(x : int366_t) return std_logic_vector is
  variable rv : std_logic_vector(365 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int366_t(x : std_logic_vector) return int366_t is
  variable rv : int366_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint367_t_to_slv(x : uint367_t) return std_logic_vector is
  variable rv : std_logic_vector(366 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint367_t(x : std_logic_vector) return uint367_t is
  variable rv : uint367_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int367_t_to_slv(x : int367_t) return std_logic_vector is
  variable rv : std_logic_vector(366 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int367_t(x : std_logic_vector) return int367_t is
  variable rv : int367_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint368_t_to_slv(x : uint368_t) return std_logic_vector is
  variable rv : std_logic_vector(367 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint368_t(x : std_logic_vector) return uint368_t is
  variable rv : uint368_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int368_t_to_slv(x : int368_t) return std_logic_vector is
  variable rv : std_logic_vector(367 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int368_t(x : std_logic_vector) return int368_t is
  variable rv : int368_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint369_t_to_slv(x : uint369_t) return std_logic_vector is
  variable rv : std_logic_vector(368 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint369_t(x : std_logic_vector) return uint369_t is
  variable rv : uint369_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int369_t_to_slv(x : int369_t) return std_logic_vector is
  variable rv : std_logic_vector(368 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int369_t(x : std_logic_vector) return int369_t is
  variable rv : int369_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint370_t_to_slv(x : uint370_t) return std_logic_vector is
  variable rv : std_logic_vector(369 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint370_t(x : std_logic_vector) return uint370_t is
  variable rv : uint370_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int370_t_to_slv(x : int370_t) return std_logic_vector is
  variable rv : std_logic_vector(369 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int370_t(x : std_logic_vector) return int370_t is
  variable rv : int370_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint371_t_to_slv(x : uint371_t) return std_logic_vector is
  variable rv : std_logic_vector(370 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint371_t(x : std_logic_vector) return uint371_t is
  variable rv : uint371_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int371_t_to_slv(x : int371_t) return std_logic_vector is
  variable rv : std_logic_vector(370 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int371_t(x : std_logic_vector) return int371_t is
  variable rv : int371_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint372_t_to_slv(x : uint372_t) return std_logic_vector is
  variable rv : std_logic_vector(371 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint372_t(x : std_logic_vector) return uint372_t is
  variable rv : uint372_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int372_t_to_slv(x : int372_t) return std_logic_vector is
  variable rv : std_logic_vector(371 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int372_t(x : std_logic_vector) return int372_t is
  variable rv : int372_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint373_t_to_slv(x : uint373_t) return std_logic_vector is
  variable rv : std_logic_vector(372 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint373_t(x : std_logic_vector) return uint373_t is
  variable rv : uint373_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int373_t_to_slv(x : int373_t) return std_logic_vector is
  variable rv : std_logic_vector(372 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int373_t(x : std_logic_vector) return int373_t is
  variable rv : int373_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint374_t_to_slv(x : uint374_t) return std_logic_vector is
  variable rv : std_logic_vector(373 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint374_t(x : std_logic_vector) return uint374_t is
  variable rv : uint374_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int374_t_to_slv(x : int374_t) return std_logic_vector is
  variable rv : std_logic_vector(373 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int374_t(x : std_logic_vector) return int374_t is
  variable rv : int374_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint375_t_to_slv(x : uint375_t) return std_logic_vector is
  variable rv : std_logic_vector(374 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint375_t(x : std_logic_vector) return uint375_t is
  variable rv : uint375_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int375_t_to_slv(x : int375_t) return std_logic_vector is
  variable rv : std_logic_vector(374 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int375_t(x : std_logic_vector) return int375_t is
  variable rv : int375_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint376_t_to_slv(x : uint376_t) return std_logic_vector is
  variable rv : std_logic_vector(375 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint376_t(x : std_logic_vector) return uint376_t is
  variable rv : uint376_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int376_t_to_slv(x : int376_t) return std_logic_vector is
  variable rv : std_logic_vector(375 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int376_t(x : std_logic_vector) return int376_t is
  variable rv : int376_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint377_t_to_slv(x : uint377_t) return std_logic_vector is
  variable rv : std_logic_vector(376 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint377_t(x : std_logic_vector) return uint377_t is
  variable rv : uint377_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int377_t_to_slv(x : int377_t) return std_logic_vector is
  variable rv : std_logic_vector(376 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int377_t(x : std_logic_vector) return int377_t is
  variable rv : int377_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint378_t_to_slv(x : uint378_t) return std_logic_vector is
  variable rv : std_logic_vector(377 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint378_t(x : std_logic_vector) return uint378_t is
  variable rv : uint378_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int378_t_to_slv(x : int378_t) return std_logic_vector is
  variable rv : std_logic_vector(377 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int378_t(x : std_logic_vector) return int378_t is
  variable rv : int378_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint379_t_to_slv(x : uint379_t) return std_logic_vector is
  variable rv : std_logic_vector(378 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint379_t(x : std_logic_vector) return uint379_t is
  variable rv : uint379_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int379_t_to_slv(x : int379_t) return std_logic_vector is
  variable rv : std_logic_vector(378 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int379_t(x : std_logic_vector) return int379_t is
  variable rv : int379_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint380_t_to_slv(x : uint380_t) return std_logic_vector is
  variable rv : std_logic_vector(379 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint380_t(x : std_logic_vector) return uint380_t is
  variable rv : uint380_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int380_t_to_slv(x : int380_t) return std_logic_vector is
  variable rv : std_logic_vector(379 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int380_t(x : std_logic_vector) return int380_t is
  variable rv : int380_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint381_t_to_slv(x : uint381_t) return std_logic_vector is
  variable rv : std_logic_vector(380 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint381_t(x : std_logic_vector) return uint381_t is
  variable rv : uint381_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int381_t_to_slv(x : int381_t) return std_logic_vector is
  variable rv : std_logic_vector(380 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int381_t(x : std_logic_vector) return int381_t is
  variable rv : int381_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint382_t_to_slv(x : uint382_t) return std_logic_vector is
  variable rv : std_logic_vector(381 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint382_t(x : std_logic_vector) return uint382_t is
  variable rv : uint382_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int382_t_to_slv(x : int382_t) return std_logic_vector is
  variable rv : std_logic_vector(381 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int382_t(x : std_logic_vector) return int382_t is
  variable rv : int382_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint383_t_to_slv(x : uint383_t) return std_logic_vector is
  variable rv : std_logic_vector(382 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint383_t(x : std_logic_vector) return uint383_t is
  variable rv : uint383_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int383_t_to_slv(x : int383_t) return std_logic_vector is
  variable rv : std_logic_vector(382 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int383_t(x : std_logic_vector) return int383_t is
  variable rv : int383_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint384_t_to_slv(x : uint384_t) return std_logic_vector is
  variable rv : std_logic_vector(383 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint384_t(x : std_logic_vector) return uint384_t is
  variable rv : uint384_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int384_t_to_slv(x : int384_t) return std_logic_vector is
  variable rv : std_logic_vector(383 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int384_t(x : std_logic_vector) return int384_t is
  variable rv : int384_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint385_t_to_slv(x : uint385_t) return std_logic_vector is
  variable rv : std_logic_vector(384 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint385_t(x : std_logic_vector) return uint385_t is
  variable rv : uint385_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int385_t_to_slv(x : int385_t) return std_logic_vector is
  variable rv : std_logic_vector(384 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int385_t(x : std_logic_vector) return int385_t is
  variable rv : int385_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint386_t_to_slv(x : uint386_t) return std_logic_vector is
  variable rv : std_logic_vector(385 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint386_t(x : std_logic_vector) return uint386_t is
  variable rv : uint386_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int386_t_to_slv(x : int386_t) return std_logic_vector is
  variable rv : std_logic_vector(385 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int386_t(x : std_logic_vector) return int386_t is
  variable rv : int386_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint387_t_to_slv(x : uint387_t) return std_logic_vector is
  variable rv : std_logic_vector(386 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint387_t(x : std_logic_vector) return uint387_t is
  variable rv : uint387_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int387_t_to_slv(x : int387_t) return std_logic_vector is
  variable rv : std_logic_vector(386 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int387_t(x : std_logic_vector) return int387_t is
  variable rv : int387_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint388_t_to_slv(x : uint388_t) return std_logic_vector is
  variable rv : std_logic_vector(387 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint388_t(x : std_logic_vector) return uint388_t is
  variable rv : uint388_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int388_t_to_slv(x : int388_t) return std_logic_vector is
  variable rv : std_logic_vector(387 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int388_t(x : std_logic_vector) return int388_t is
  variable rv : int388_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint389_t_to_slv(x : uint389_t) return std_logic_vector is
  variable rv : std_logic_vector(388 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint389_t(x : std_logic_vector) return uint389_t is
  variable rv : uint389_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int389_t_to_slv(x : int389_t) return std_logic_vector is
  variable rv : std_logic_vector(388 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int389_t(x : std_logic_vector) return int389_t is
  variable rv : int389_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint390_t_to_slv(x : uint390_t) return std_logic_vector is
  variable rv : std_logic_vector(389 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint390_t(x : std_logic_vector) return uint390_t is
  variable rv : uint390_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int390_t_to_slv(x : int390_t) return std_logic_vector is
  variable rv : std_logic_vector(389 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int390_t(x : std_logic_vector) return int390_t is
  variable rv : int390_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint391_t_to_slv(x : uint391_t) return std_logic_vector is
  variable rv : std_logic_vector(390 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint391_t(x : std_logic_vector) return uint391_t is
  variable rv : uint391_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int391_t_to_slv(x : int391_t) return std_logic_vector is
  variable rv : std_logic_vector(390 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int391_t(x : std_logic_vector) return int391_t is
  variable rv : int391_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint392_t_to_slv(x : uint392_t) return std_logic_vector is
  variable rv : std_logic_vector(391 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint392_t(x : std_logic_vector) return uint392_t is
  variable rv : uint392_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int392_t_to_slv(x : int392_t) return std_logic_vector is
  variable rv : std_logic_vector(391 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int392_t(x : std_logic_vector) return int392_t is
  variable rv : int392_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint393_t_to_slv(x : uint393_t) return std_logic_vector is
  variable rv : std_logic_vector(392 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint393_t(x : std_logic_vector) return uint393_t is
  variable rv : uint393_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int393_t_to_slv(x : int393_t) return std_logic_vector is
  variable rv : std_logic_vector(392 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int393_t(x : std_logic_vector) return int393_t is
  variable rv : int393_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint394_t_to_slv(x : uint394_t) return std_logic_vector is
  variable rv : std_logic_vector(393 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint394_t(x : std_logic_vector) return uint394_t is
  variable rv : uint394_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int394_t_to_slv(x : int394_t) return std_logic_vector is
  variable rv : std_logic_vector(393 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int394_t(x : std_logic_vector) return int394_t is
  variable rv : int394_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint395_t_to_slv(x : uint395_t) return std_logic_vector is
  variable rv : std_logic_vector(394 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint395_t(x : std_logic_vector) return uint395_t is
  variable rv : uint395_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int395_t_to_slv(x : int395_t) return std_logic_vector is
  variable rv : std_logic_vector(394 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int395_t(x : std_logic_vector) return int395_t is
  variable rv : int395_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint396_t_to_slv(x : uint396_t) return std_logic_vector is
  variable rv : std_logic_vector(395 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint396_t(x : std_logic_vector) return uint396_t is
  variable rv : uint396_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int396_t_to_slv(x : int396_t) return std_logic_vector is
  variable rv : std_logic_vector(395 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int396_t(x : std_logic_vector) return int396_t is
  variable rv : int396_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint397_t_to_slv(x : uint397_t) return std_logic_vector is
  variable rv : std_logic_vector(396 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint397_t(x : std_logic_vector) return uint397_t is
  variable rv : uint397_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int397_t_to_slv(x : int397_t) return std_logic_vector is
  variable rv : std_logic_vector(396 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int397_t(x : std_logic_vector) return int397_t is
  variable rv : int397_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint398_t_to_slv(x : uint398_t) return std_logic_vector is
  variable rv : std_logic_vector(397 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint398_t(x : std_logic_vector) return uint398_t is
  variable rv : uint398_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int398_t_to_slv(x : int398_t) return std_logic_vector is
  variable rv : std_logic_vector(397 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int398_t(x : std_logic_vector) return int398_t is
  variable rv : int398_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint399_t_to_slv(x : uint399_t) return std_logic_vector is
  variable rv : std_logic_vector(398 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint399_t(x : std_logic_vector) return uint399_t is
  variable rv : uint399_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int399_t_to_slv(x : int399_t) return std_logic_vector is
  variable rv : std_logic_vector(398 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int399_t(x : std_logic_vector) return int399_t is
  variable rv : int399_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint400_t_to_slv(x : uint400_t) return std_logic_vector is
  variable rv : std_logic_vector(399 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint400_t(x : std_logic_vector) return uint400_t is
  variable rv : uint400_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int400_t_to_slv(x : int400_t) return std_logic_vector is
  variable rv : std_logic_vector(399 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int400_t(x : std_logic_vector) return int400_t is
  variable rv : int400_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint401_t_to_slv(x : uint401_t) return std_logic_vector is
  variable rv : std_logic_vector(400 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint401_t(x : std_logic_vector) return uint401_t is
  variable rv : uint401_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int401_t_to_slv(x : int401_t) return std_logic_vector is
  variable rv : std_logic_vector(400 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int401_t(x : std_logic_vector) return int401_t is
  variable rv : int401_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint402_t_to_slv(x : uint402_t) return std_logic_vector is
  variable rv : std_logic_vector(401 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint402_t(x : std_logic_vector) return uint402_t is
  variable rv : uint402_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int402_t_to_slv(x : int402_t) return std_logic_vector is
  variable rv : std_logic_vector(401 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int402_t(x : std_logic_vector) return int402_t is
  variable rv : int402_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint403_t_to_slv(x : uint403_t) return std_logic_vector is
  variable rv : std_logic_vector(402 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint403_t(x : std_logic_vector) return uint403_t is
  variable rv : uint403_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int403_t_to_slv(x : int403_t) return std_logic_vector is
  variable rv : std_logic_vector(402 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int403_t(x : std_logic_vector) return int403_t is
  variable rv : int403_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint404_t_to_slv(x : uint404_t) return std_logic_vector is
  variable rv : std_logic_vector(403 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint404_t(x : std_logic_vector) return uint404_t is
  variable rv : uint404_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int404_t_to_slv(x : int404_t) return std_logic_vector is
  variable rv : std_logic_vector(403 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int404_t(x : std_logic_vector) return int404_t is
  variable rv : int404_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint405_t_to_slv(x : uint405_t) return std_logic_vector is
  variable rv : std_logic_vector(404 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint405_t(x : std_logic_vector) return uint405_t is
  variable rv : uint405_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int405_t_to_slv(x : int405_t) return std_logic_vector is
  variable rv : std_logic_vector(404 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int405_t(x : std_logic_vector) return int405_t is
  variable rv : int405_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint406_t_to_slv(x : uint406_t) return std_logic_vector is
  variable rv : std_logic_vector(405 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint406_t(x : std_logic_vector) return uint406_t is
  variable rv : uint406_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int406_t_to_slv(x : int406_t) return std_logic_vector is
  variable rv : std_logic_vector(405 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int406_t(x : std_logic_vector) return int406_t is
  variable rv : int406_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint407_t_to_slv(x : uint407_t) return std_logic_vector is
  variable rv : std_logic_vector(406 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint407_t(x : std_logic_vector) return uint407_t is
  variable rv : uint407_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int407_t_to_slv(x : int407_t) return std_logic_vector is
  variable rv : std_logic_vector(406 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int407_t(x : std_logic_vector) return int407_t is
  variable rv : int407_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint408_t_to_slv(x : uint408_t) return std_logic_vector is
  variable rv : std_logic_vector(407 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint408_t(x : std_logic_vector) return uint408_t is
  variable rv : uint408_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int408_t_to_slv(x : int408_t) return std_logic_vector is
  variable rv : std_logic_vector(407 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int408_t(x : std_logic_vector) return int408_t is
  variable rv : int408_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint409_t_to_slv(x : uint409_t) return std_logic_vector is
  variable rv : std_logic_vector(408 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint409_t(x : std_logic_vector) return uint409_t is
  variable rv : uint409_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int409_t_to_slv(x : int409_t) return std_logic_vector is
  variable rv : std_logic_vector(408 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int409_t(x : std_logic_vector) return int409_t is
  variable rv : int409_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint410_t_to_slv(x : uint410_t) return std_logic_vector is
  variable rv : std_logic_vector(409 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint410_t(x : std_logic_vector) return uint410_t is
  variable rv : uint410_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int410_t_to_slv(x : int410_t) return std_logic_vector is
  variable rv : std_logic_vector(409 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int410_t(x : std_logic_vector) return int410_t is
  variable rv : int410_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint411_t_to_slv(x : uint411_t) return std_logic_vector is
  variable rv : std_logic_vector(410 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint411_t(x : std_logic_vector) return uint411_t is
  variable rv : uint411_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int411_t_to_slv(x : int411_t) return std_logic_vector is
  variable rv : std_logic_vector(410 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int411_t(x : std_logic_vector) return int411_t is
  variable rv : int411_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint412_t_to_slv(x : uint412_t) return std_logic_vector is
  variable rv : std_logic_vector(411 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint412_t(x : std_logic_vector) return uint412_t is
  variable rv : uint412_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int412_t_to_slv(x : int412_t) return std_logic_vector is
  variable rv : std_logic_vector(411 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int412_t(x : std_logic_vector) return int412_t is
  variable rv : int412_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint413_t_to_slv(x : uint413_t) return std_logic_vector is
  variable rv : std_logic_vector(412 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint413_t(x : std_logic_vector) return uint413_t is
  variable rv : uint413_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int413_t_to_slv(x : int413_t) return std_logic_vector is
  variable rv : std_logic_vector(412 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int413_t(x : std_logic_vector) return int413_t is
  variable rv : int413_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint414_t_to_slv(x : uint414_t) return std_logic_vector is
  variable rv : std_logic_vector(413 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint414_t(x : std_logic_vector) return uint414_t is
  variable rv : uint414_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int414_t_to_slv(x : int414_t) return std_logic_vector is
  variable rv : std_logic_vector(413 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int414_t(x : std_logic_vector) return int414_t is
  variable rv : int414_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint415_t_to_slv(x : uint415_t) return std_logic_vector is
  variable rv : std_logic_vector(414 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint415_t(x : std_logic_vector) return uint415_t is
  variable rv : uint415_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int415_t_to_slv(x : int415_t) return std_logic_vector is
  variable rv : std_logic_vector(414 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int415_t(x : std_logic_vector) return int415_t is
  variable rv : int415_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint416_t_to_slv(x : uint416_t) return std_logic_vector is
  variable rv : std_logic_vector(415 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint416_t(x : std_logic_vector) return uint416_t is
  variable rv : uint416_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int416_t_to_slv(x : int416_t) return std_logic_vector is
  variable rv : std_logic_vector(415 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int416_t(x : std_logic_vector) return int416_t is
  variable rv : int416_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint417_t_to_slv(x : uint417_t) return std_logic_vector is
  variable rv : std_logic_vector(416 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint417_t(x : std_logic_vector) return uint417_t is
  variable rv : uint417_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int417_t_to_slv(x : int417_t) return std_logic_vector is
  variable rv : std_logic_vector(416 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int417_t(x : std_logic_vector) return int417_t is
  variable rv : int417_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint418_t_to_slv(x : uint418_t) return std_logic_vector is
  variable rv : std_logic_vector(417 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint418_t(x : std_logic_vector) return uint418_t is
  variable rv : uint418_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int418_t_to_slv(x : int418_t) return std_logic_vector is
  variable rv : std_logic_vector(417 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int418_t(x : std_logic_vector) return int418_t is
  variable rv : int418_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint419_t_to_slv(x : uint419_t) return std_logic_vector is
  variable rv : std_logic_vector(418 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint419_t(x : std_logic_vector) return uint419_t is
  variable rv : uint419_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int419_t_to_slv(x : int419_t) return std_logic_vector is
  variable rv : std_logic_vector(418 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int419_t(x : std_logic_vector) return int419_t is
  variable rv : int419_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint420_t_to_slv(x : uint420_t) return std_logic_vector is
  variable rv : std_logic_vector(419 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint420_t(x : std_logic_vector) return uint420_t is
  variable rv : uint420_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int420_t_to_slv(x : int420_t) return std_logic_vector is
  variable rv : std_logic_vector(419 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int420_t(x : std_logic_vector) return int420_t is
  variable rv : int420_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint421_t_to_slv(x : uint421_t) return std_logic_vector is
  variable rv : std_logic_vector(420 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint421_t(x : std_logic_vector) return uint421_t is
  variable rv : uint421_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int421_t_to_slv(x : int421_t) return std_logic_vector is
  variable rv : std_logic_vector(420 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int421_t(x : std_logic_vector) return int421_t is
  variable rv : int421_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint422_t_to_slv(x : uint422_t) return std_logic_vector is
  variable rv : std_logic_vector(421 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint422_t(x : std_logic_vector) return uint422_t is
  variable rv : uint422_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int422_t_to_slv(x : int422_t) return std_logic_vector is
  variable rv : std_logic_vector(421 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int422_t(x : std_logic_vector) return int422_t is
  variable rv : int422_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint423_t_to_slv(x : uint423_t) return std_logic_vector is
  variable rv : std_logic_vector(422 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint423_t(x : std_logic_vector) return uint423_t is
  variable rv : uint423_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int423_t_to_slv(x : int423_t) return std_logic_vector is
  variable rv : std_logic_vector(422 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int423_t(x : std_logic_vector) return int423_t is
  variable rv : int423_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint424_t_to_slv(x : uint424_t) return std_logic_vector is
  variable rv : std_logic_vector(423 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint424_t(x : std_logic_vector) return uint424_t is
  variable rv : uint424_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int424_t_to_slv(x : int424_t) return std_logic_vector is
  variable rv : std_logic_vector(423 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int424_t(x : std_logic_vector) return int424_t is
  variable rv : int424_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint425_t_to_slv(x : uint425_t) return std_logic_vector is
  variable rv : std_logic_vector(424 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint425_t(x : std_logic_vector) return uint425_t is
  variable rv : uint425_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int425_t_to_slv(x : int425_t) return std_logic_vector is
  variable rv : std_logic_vector(424 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int425_t(x : std_logic_vector) return int425_t is
  variable rv : int425_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint426_t_to_slv(x : uint426_t) return std_logic_vector is
  variable rv : std_logic_vector(425 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint426_t(x : std_logic_vector) return uint426_t is
  variable rv : uint426_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int426_t_to_slv(x : int426_t) return std_logic_vector is
  variable rv : std_logic_vector(425 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int426_t(x : std_logic_vector) return int426_t is
  variable rv : int426_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint427_t_to_slv(x : uint427_t) return std_logic_vector is
  variable rv : std_logic_vector(426 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint427_t(x : std_logic_vector) return uint427_t is
  variable rv : uint427_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int427_t_to_slv(x : int427_t) return std_logic_vector is
  variable rv : std_logic_vector(426 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int427_t(x : std_logic_vector) return int427_t is
  variable rv : int427_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint428_t_to_slv(x : uint428_t) return std_logic_vector is
  variable rv : std_logic_vector(427 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint428_t(x : std_logic_vector) return uint428_t is
  variable rv : uint428_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int428_t_to_slv(x : int428_t) return std_logic_vector is
  variable rv : std_logic_vector(427 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int428_t(x : std_logic_vector) return int428_t is
  variable rv : int428_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint429_t_to_slv(x : uint429_t) return std_logic_vector is
  variable rv : std_logic_vector(428 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint429_t(x : std_logic_vector) return uint429_t is
  variable rv : uint429_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int429_t_to_slv(x : int429_t) return std_logic_vector is
  variable rv : std_logic_vector(428 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int429_t(x : std_logic_vector) return int429_t is
  variable rv : int429_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint430_t_to_slv(x : uint430_t) return std_logic_vector is
  variable rv : std_logic_vector(429 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint430_t(x : std_logic_vector) return uint430_t is
  variable rv : uint430_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int430_t_to_slv(x : int430_t) return std_logic_vector is
  variable rv : std_logic_vector(429 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int430_t(x : std_logic_vector) return int430_t is
  variable rv : int430_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint431_t_to_slv(x : uint431_t) return std_logic_vector is
  variable rv : std_logic_vector(430 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint431_t(x : std_logic_vector) return uint431_t is
  variable rv : uint431_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int431_t_to_slv(x : int431_t) return std_logic_vector is
  variable rv : std_logic_vector(430 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int431_t(x : std_logic_vector) return int431_t is
  variable rv : int431_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint432_t_to_slv(x : uint432_t) return std_logic_vector is
  variable rv : std_logic_vector(431 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint432_t(x : std_logic_vector) return uint432_t is
  variable rv : uint432_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int432_t_to_slv(x : int432_t) return std_logic_vector is
  variable rv : std_logic_vector(431 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int432_t(x : std_logic_vector) return int432_t is
  variable rv : int432_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint433_t_to_slv(x : uint433_t) return std_logic_vector is
  variable rv : std_logic_vector(432 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint433_t(x : std_logic_vector) return uint433_t is
  variable rv : uint433_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int433_t_to_slv(x : int433_t) return std_logic_vector is
  variable rv : std_logic_vector(432 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int433_t(x : std_logic_vector) return int433_t is
  variable rv : int433_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint434_t_to_slv(x : uint434_t) return std_logic_vector is
  variable rv : std_logic_vector(433 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint434_t(x : std_logic_vector) return uint434_t is
  variable rv : uint434_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int434_t_to_slv(x : int434_t) return std_logic_vector is
  variable rv : std_logic_vector(433 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int434_t(x : std_logic_vector) return int434_t is
  variable rv : int434_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint435_t_to_slv(x : uint435_t) return std_logic_vector is
  variable rv : std_logic_vector(434 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint435_t(x : std_logic_vector) return uint435_t is
  variable rv : uint435_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int435_t_to_slv(x : int435_t) return std_logic_vector is
  variable rv : std_logic_vector(434 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int435_t(x : std_logic_vector) return int435_t is
  variable rv : int435_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint436_t_to_slv(x : uint436_t) return std_logic_vector is
  variable rv : std_logic_vector(435 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint436_t(x : std_logic_vector) return uint436_t is
  variable rv : uint436_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int436_t_to_slv(x : int436_t) return std_logic_vector is
  variable rv : std_logic_vector(435 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int436_t(x : std_logic_vector) return int436_t is
  variable rv : int436_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint437_t_to_slv(x : uint437_t) return std_logic_vector is
  variable rv : std_logic_vector(436 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint437_t(x : std_logic_vector) return uint437_t is
  variable rv : uint437_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int437_t_to_slv(x : int437_t) return std_logic_vector is
  variable rv : std_logic_vector(436 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int437_t(x : std_logic_vector) return int437_t is
  variable rv : int437_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint438_t_to_slv(x : uint438_t) return std_logic_vector is
  variable rv : std_logic_vector(437 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint438_t(x : std_logic_vector) return uint438_t is
  variable rv : uint438_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int438_t_to_slv(x : int438_t) return std_logic_vector is
  variable rv : std_logic_vector(437 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int438_t(x : std_logic_vector) return int438_t is
  variable rv : int438_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint439_t_to_slv(x : uint439_t) return std_logic_vector is
  variable rv : std_logic_vector(438 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint439_t(x : std_logic_vector) return uint439_t is
  variable rv : uint439_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int439_t_to_slv(x : int439_t) return std_logic_vector is
  variable rv : std_logic_vector(438 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int439_t(x : std_logic_vector) return int439_t is
  variable rv : int439_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint440_t_to_slv(x : uint440_t) return std_logic_vector is
  variable rv : std_logic_vector(439 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint440_t(x : std_logic_vector) return uint440_t is
  variable rv : uint440_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int440_t_to_slv(x : int440_t) return std_logic_vector is
  variable rv : std_logic_vector(439 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int440_t(x : std_logic_vector) return int440_t is
  variable rv : int440_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint441_t_to_slv(x : uint441_t) return std_logic_vector is
  variable rv : std_logic_vector(440 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint441_t(x : std_logic_vector) return uint441_t is
  variable rv : uint441_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int441_t_to_slv(x : int441_t) return std_logic_vector is
  variable rv : std_logic_vector(440 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int441_t(x : std_logic_vector) return int441_t is
  variable rv : int441_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint442_t_to_slv(x : uint442_t) return std_logic_vector is
  variable rv : std_logic_vector(441 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint442_t(x : std_logic_vector) return uint442_t is
  variable rv : uint442_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int442_t_to_slv(x : int442_t) return std_logic_vector is
  variable rv : std_logic_vector(441 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int442_t(x : std_logic_vector) return int442_t is
  variable rv : int442_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint443_t_to_slv(x : uint443_t) return std_logic_vector is
  variable rv : std_logic_vector(442 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint443_t(x : std_logic_vector) return uint443_t is
  variable rv : uint443_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int443_t_to_slv(x : int443_t) return std_logic_vector is
  variable rv : std_logic_vector(442 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int443_t(x : std_logic_vector) return int443_t is
  variable rv : int443_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint444_t_to_slv(x : uint444_t) return std_logic_vector is
  variable rv : std_logic_vector(443 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint444_t(x : std_logic_vector) return uint444_t is
  variable rv : uint444_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int444_t_to_slv(x : int444_t) return std_logic_vector is
  variable rv : std_logic_vector(443 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int444_t(x : std_logic_vector) return int444_t is
  variable rv : int444_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint445_t_to_slv(x : uint445_t) return std_logic_vector is
  variable rv : std_logic_vector(444 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint445_t(x : std_logic_vector) return uint445_t is
  variable rv : uint445_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int445_t_to_slv(x : int445_t) return std_logic_vector is
  variable rv : std_logic_vector(444 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int445_t(x : std_logic_vector) return int445_t is
  variable rv : int445_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint446_t_to_slv(x : uint446_t) return std_logic_vector is
  variable rv : std_logic_vector(445 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint446_t(x : std_logic_vector) return uint446_t is
  variable rv : uint446_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int446_t_to_slv(x : int446_t) return std_logic_vector is
  variable rv : std_logic_vector(445 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int446_t(x : std_logic_vector) return int446_t is
  variable rv : int446_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint447_t_to_slv(x : uint447_t) return std_logic_vector is
  variable rv : std_logic_vector(446 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint447_t(x : std_logic_vector) return uint447_t is
  variable rv : uint447_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int447_t_to_slv(x : int447_t) return std_logic_vector is
  variable rv : std_logic_vector(446 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int447_t(x : std_logic_vector) return int447_t is
  variable rv : int447_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint448_t_to_slv(x : uint448_t) return std_logic_vector is
  variable rv : std_logic_vector(447 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint448_t(x : std_logic_vector) return uint448_t is
  variable rv : uint448_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int448_t_to_slv(x : int448_t) return std_logic_vector is
  variable rv : std_logic_vector(447 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int448_t(x : std_logic_vector) return int448_t is
  variable rv : int448_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint449_t_to_slv(x : uint449_t) return std_logic_vector is
  variable rv : std_logic_vector(448 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint449_t(x : std_logic_vector) return uint449_t is
  variable rv : uint449_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int449_t_to_slv(x : int449_t) return std_logic_vector is
  variable rv : std_logic_vector(448 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int449_t(x : std_logic_vector) return int449_t is
  variable rv : int449_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint450_t_to_slv(x : uint450_t) return std_logic_vector is
  variable rv : std_logic_vector(449 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint450_t(x : std_logic_vector) return uint450_t is
  variable rv : uint450_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int450_t_to_slv(x : int450_t) return std_logic_vector is
  variable rv : std_logic_vector(449 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int450_t(x : std_logic_vector) return int450_t is
  variable rv : int450_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint451_t_to_slv(x : uint451_t) return std_logic_vector is
  variable rv : std_logic_vector(450 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint451_t(x : std_logic_vector) return uint451_t is
  variable rv : uint451_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int451_t_to_slv(x : int451_t) return std_logic_vector is
  variable rv : std_logic_vector(450 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int451_t(x : std_logic_vector) return int451_t is
  variable rv : int451_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint452_t_to_slv(x : uint452_t) return std_logic_vector is
  variable rv : std_logic_vector(451 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint452_t(x : std_logic_vector) return uint452_t is
  variable rv : uint452_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int452_t_to_slv(x : int452_t) return std_logic_vector is
  variable rv : std_logic_vector(451 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int452_t(x : std_logic_vector) return int452_t is
  variable rv : int452_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint453_t_to_slv(x : uint453_t) return std_logic_vector is
  variable rv : std_logic_vector(452 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint453_t(x : std_logic_vector) return uint453_t is
  variable rv : uint453_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int453_t_to_slv(x : int453_t) return std_logic_vector is
  variable rv : std_logic_vector(452 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int453_t(x : std_logic_vector) return int453_t is
  variable rv : int453_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint454_t_to_slv(x : uint454_t) return std_logic_vector is
  variable rv : std_logic_vector(453 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint454_t(x : std_logic_vector) return uint454_t is
  variable rv : uint454_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int454_t_to_slv(x : int454_t) return std_logic_vector is
  variable rv : std_logic_vector(453 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int454_t(x : std_logic_vector) return int454_t is
  variable rv : int454_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint455_t_to_slv(x : uint455_t) return std_logic_vector is
  variable rv : std_logic_vector(454 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint455_t(x : std_logic_vector) return uint455_t is
  variable rv : uint455_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int455_t_to_slv(x : int455_t) return std_logic_vector is
  variable rv : std_logic_vector(454 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int455_t(x : std_logic_vector) return int455_t is
  variable rv : int455_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint456_t_to_slv(x : uint456_t) return std_logic_vector is
  variable rv : std_logic_vector(455 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint456_t(x : std_logic_vector) return uint456_t is
  variable rv : uint456_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int456_t_to_slv(x : int456_t) return std_logic_vector is
  variable rv : std_logic_vector(455 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int456_t(x : std_logic_vector) return int456_t is
  variable rv : int456_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint457_t_to_slv(x : uint457_t) return std_logic_vector is
  variable rv : std_logic_vector(456 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint457_t(x : std_logic_vector) return uint457_t is
  variable rv : uint457_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int457_t_to_slv(x : int457_t) return std_logic_vector is
  variable rv : std_logic_vector(456 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int457_t(x : std_logic_vector) return int457_t is
  variable rv : int457_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint458_t_to_slv(x : uint458_t) return std_logic_vector is
  variable rv : std_logic_vector(457 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint458_t(x : std_logic_vector) return uint458_t is
  variable rv : uint458_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int458_t_to_slv(x : int458_t) return std_logic_vector is
  variable rv : std_logic_vector(457 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int458_t(x : std_logic_vector) return int458_t is
  variable rv : int458_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint459_t_to_slv(x : uint459_t) return std_logic_vector is
  variable rv : std_logic_vector(458 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint459_t(x : std_logic_vector) return uint459_t is
  variable rv : uint459_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int459_t_to_slv(x : int459_t) return std_logic_vector is
  variable rv : std_logic_vector(458 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int459_t(x : std_logic_vector) return int459_t is
  variable rv : int459_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint460_t_to_slv(x : uint460_t) return std_logic_vector is
  variable rv : std_logic_vector(459 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint460_t(x : std_logic_vector) return uint460_t is
  variable rv : uint460_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int460_t_to_slv(x : int460_t) return std_logic_vector is
  variable rv : std_logic_vector(459 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int460_t(x : std_logic_vector) return int460_t is
  variable rv : int460_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint461_t_to_slv(x : uint461_t) return std_logic_vector is
  variable rv : std_logic_vector(460 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint461_t(x : std_logic_vector) return uint461_t is
  variable rv : uint461_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int461_t_to_slv(x : int461_t) return std_logic_vector is
  variable rv : std_logic_vector(460 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int461_t(x : std_logic_vector) return int461_t is
  variable rv : int461_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint462_t_to_slv(x : uint462_t) return std_logic_vector is
  variable rv : std_logic_vector(461 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint462_t(x : std_logic_vector) return uint462_t is
  variable rv : uint462_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int462_t_to_slv(x : int462_t) return std_logic_vector is
  variable rv : std_logic_vector(461 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int462_t(x : std_logic_vector) return int462_t is
  variable rv : int462_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint463_t_to_slv(x : uint463_t) return std_logic_vector is
  variable rv : std_logic_vector(462 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint463_t(x : std_logic_vector) return uint463_t is
  variable rv : uint463_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int463_t_to_slv(x : int463_t) return std_logic_vector is
  variable rv : std_logic_vector(462 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int463_t(x : std_logic_vector) return int463_t is
  variable rv : int463_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint464_t_to_slv(x : uint464_t) return std_logic_vector is
  variable rv : std_logic_vector(463 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint464_t(x : std_logic_vector) return uint464_t is
  variable rv : uint464_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int464_t_to_slv(x : int464_t) return std_logic_vector is
  variable rv : std_logic_vector(463 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int464_t(x : std_logic_vector) return int464_t is
  variable rv : int464_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint465_t_to_slv(x : uint465_t) return std_logic_vector is
  variable rv : std_logic_vector(464 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint465_t(x : std_logic_vector) return uint465_t is
  variable rv : uint465_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int465_t_to_slv(x : int465_t) return std_logic_vector is
  variable rv : std_logic_vector(464 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int465_t(x : std_logic_vector) return int465_t is
  variable rv : int465_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint466_t_to_slv(x : uint466_t) return std_logic_vector is
  variable rv : std_logic_vector(465 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint466_t(x : std_logic_vector) return uint466_t is
  variable rv : uint466_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int466_t_to_slv(x : int466_t) return std_logic_vector is
  variable rv : std_logic_vector(465 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int466_t(x : std_logic_vector) return int466_t is
  variable rv : int466_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint467_t_to_slv(x : uint467_t) return std_logic_vector is
  variable rv : std_logic_vector(466 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint467_t(x : std_logic_vector) return uint467_t is
  variable rv : uint467_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int467_t_to_slv(x : int467_t) return std_logic_vector is
  variable rv : std_logic_vector(466 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int467_t(x : std_logic_vector) return int467_t is
  variable rv : int467_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint468_t_to_slv(x : uint468_t) return std_logic_vector is
  variable rv : std_logic_vector(467 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint468_t(x : std_logic_vector) return uint468_t is
  variable rv : uint468_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int468_t_to_slv(x : int468_t) return std_logic_vector is
  variable rv : std_logic_vector(467 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int468_t(x : std_logic_vector) return int468_t is
  variable rv : int468_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint469_t_to_slv(x : uint469_t) return std_logic_vector is
  variable rv : std_logic_vector(468 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint469_t(x : std_logic_vector) return uint469_t is
  variable rv : uint469_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int469_t_to_slv(x : int469_t) return std_logic_vector is
  variable rv : std_logic_vector(468 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int469_t(x : std_logic_vector) return int469_t is
  variable rv : int469_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint470_t_to_slv(x : uint470_t) return std_logic_vector is
  variable rv : std_logic_vector(469 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint470_t(x : std_logic_vector) return uint470_t is
  variable rv : uint470_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int470_t_to_slv(x : int470_t) return std_logic_vector is
  variable rv : std_logic_vector(469 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int470_t(x : std_logic_vector) return int470_t is
  variable rv : int470_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint471_t_to_slv(x : uint471_t) return std_logic_vector is
  variable rv : std_logic_vector(470 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint471_t(x : std_logic_vector) return uint471_t is
  variable rv : uint471_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int471_t_to_slv(x : int471_t) return std_logic_vector is
  variable rv : std_logic_vector(470 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int471_t(x : std_logic_vector) return int471_t is
  variable rv : int471_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint472_t_to_slv(x : uint472_t) return std_logic_vector is
  variable rv : std_logic_vector(471 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint472_t(x : std_logic_vector) return uint472_t is
  variable rv : uint472_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int472_t_to_slv(x : int472_t) return std_logic_vector is
  variable rv : std_logic_vector(471 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int472_t(x : std_logic_vector) return int472_t is
  variable rv : int472_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint473_t_to_slv(x : uint473_t) return std_logic_vector is
  variable rv : std_logic_vector(472 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint473_t(x : std_logic_vector) return uint473_t is
  variable rv : uint473_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int473_t_to_slv(x : int473_t) return std_logic_vector is
  variable rv : std_logic_vector(472 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int473_t(x : std_logic_vector) return int473_t is
  variable rv : int473_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint474_t_to_slv(x : uint474_t) return std_logic_vector is
  variable rv : std_logic_vector(473 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint474_t(x : std_logic_vector) return uint474_t is
  variable rv : uint474_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int474_t_to_slv(x : int474_t) return std_logic_vector is
  variable rv : std_logic_vector(473 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int474_t(x : std_logic_vector) return int474_t is
  variable rv : int474_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint475_t_to_slv(x : uint475_t) return std_logic_vector is
  variable rv : std_logic_vector(474 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint475_t(x : std_logic_vector) return uint475_t is
  variable rv : uint475_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int475_t_to_slv(x : int475_t) return std_logic_vector is
  variable rv : std_logic_vector(474 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int475_t(x : std_logic_vector) return int475_t is
  variable rv : int475_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint476_t_to_slv(x : uint476_t) return std_logic_vector is
  variable rv : std_logic_vector(475 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint476_t(x : std_logic_vector) return uint476_t is
  variable rv : uint476_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int476_t_to_slv(x : int476_t) return std_logic_vector is
  variable rv : std_logic_vector(475 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int476_t(x : std_logic_vector) return int476_t is
  variable rv : int476_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint477_t_to_slv(x : uint477_t) return std_logic_vector is
  variable rv : std_logic_vector(476 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint477_t(x : std_logic_vector) return uint477_t is
  variable rv : uint477_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int477_t_to_slv(x : int477_t) return std_logic_vector is
  variable rv : std_logic_vector(476 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int477_t(x : std_logic_vector) return int477_t is
  variable rv : int477_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint478_t_to_slv(x : uint478_t) return std_logic_vector is
  variable rv : std_logic_vector(477 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint478_t(x : std_logic_vector) return uint478_t is
  variable rv : uint478_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int478_t_to_slv(x : int478_t) return std_logic_vector is
  variable rv : std_logic_vector(477 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int478_t(x : std_logic_vector) return int478_t is
  variable rv : int478_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint479_t_to_slv(x : uint479_t) return std_logic_vector is
  variable rv : std_logic_vector(478 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint479_t(x : std_logic_vector) return uint479_t is
  variable rv : uint479_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int479_t_to_slv(x : int479_t) return std_logic_vector is
  variable rv : std_logic_vector(478 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int479_t(x : std_logic_vector) return int479_t is
  variable rv : int479_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint480_t_to_slv(x : uint480_t) return std_logic_vector is
  variable rv : std_logic_vector(479 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint480_t(x : std_logic_vector) return uint480_t is
  variable rv : uint480_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int480_t_to_slv(x : int480_t) return std_logic_vector is
  variable rv : std_logic_vector(479 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int480_t(x : std_logic_vector) return int480_t is
  variable rv : int480_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint481_t_to_slv(x : uint481_t) return std_logic_vector is
  variable rv : std_logic_vector(480 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint481_t(x : std_logic_vector) return uint481_t is
  variable rv : uint481_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int481_t_to_slv(x : int481_t) return std_logic_vector is
  variable rv : std_logic_vector(480 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int481_t(x : std_logic_vector) return int481_t is
  variable rv : int481_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint482_t_to_slv(x : uint482_t) return std_logic_vector is
  variable rv : std_logic_vector(481 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint482_t(x : std_logic_vector) return uint482_t is
  variable rv : uint482_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int482_t_to_slv(x : int482_t) return std_logic_vector is
  variable rv : std_logic_vector(481 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int482_t(x : std_logic_vector) return int482_t is
  variable rv : int482_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint483_t_to_slv(x : uint483_t) return std_logic_vector is
  variable rv : std_logic_vector(482 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint483_t(x : std_logic_vector) return uint483_t is
  variable rv : uint483_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int483_t_to_slv(x : int483_t) return std_logic_vector is
  variable rv : std_logic_vector(482 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int483_t(x : std_logic_vector) return int483_t is
  variable rv : int483_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint484_t_to_slv(x : uint484_t) return std_logic_vector is
  variable rv : std_logic_vector(483 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint484_t(x : std_logic_vector) return uint484_t is
  variable rv : uint484_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int484_t_to_slv(x : int484_t) return std_logic_vector is
  variable rv : std_logic_vector(483 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int484_t(x : std_logic_vector) return int484_t is
  variable rv : int484_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint485_t_to_slv(x : uint485_t) return std_logic_vector is
  variable rv : std_logic_vector(484 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint485_t(x : std_logic_vector) return uint485_t is
  variable rv : uint485_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int485_t_to_slv(x : int485_t) return std_logic_vector is
  variable rv : std_logic_vector(484 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int485_t(x : std_logic_vector) return int485_t is
  variable rv : int485_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint486_t_to_slv(x : uint486_t) return std_logic_vector is
  variable rv : std_logic_vector(485 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint486_t(x : std_logic_vector) return uint486_t is
  variable rv : uint486_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int486_t_to_slv(x : int486_t) return std_logic_vector is
  variable rv : std_logic_vector(485 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int486_t(x : std_logic_vector) return int486_t is
  variable rv : int486_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint487_t_to_slv(x : uint487_t) return std_logic_vector is
  variable rv : std_logic_vector(486 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint487_t(x : std_logic_vector) return uint487_t is
  variable rv : uint487_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int487_t_to_slv(x : int487_t) return std_logic_vector is
  variable rv : std_logic_vector(486 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int487_t(x : std_logic_vector) return int487_t is
  variable rv : int487_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint488_t_to_slv(x : uint488_t) return std_logic_vector is
  variable rv : std_logic_vector(487 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint488_t(x : std_logic_vector) return uint488_t is
  variable rv : uint488_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int488_t_to_slv(x : int488_t) return std_logic_vector is
  variable rv : std_logic_vector(487 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int488_t(x : std_logic_vector) return int488_t is
  variable rv : int488_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint489_t_to_slv(x : uint489_t) return std_logic_vector is
  variable rv : std_logic_vector(488 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint489_t(x : std_logic_vector) return uint489_t is
  variable rv : uint489_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int489_t_to_slv(x : int489_t) return std_logic_vector is
  variable rv : std_logic_vector(488 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int489_t(x : std_logic_vector) return int489_t is
  variable rv : int489_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint490_t_to_slv(x : uint490_t) return std_logic_vector is
  variable rv : std_logic_vector(489 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint490_t(x : std_logic_vector) return uint490_t is
  variable rv : uint490_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int490_t_to_slv(x : int490_t) return std_logic_vector is
  variable rv : std_logic_vector(489 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int490_t(x : std_logic_vector) return int490_t is
  variable rv : int490_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint491_t_to_slv(x : uint491_t) return std_logic_vector is
  variable rv : std_logic_vector(490 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint491_t(x : std_logic_vector) return uint491_t is
  variable rv : uint491_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int491_t_to_slv(x : int491_t) return std_logic_vector is
  variable rv : std_logic_vector(490 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int491_t(x : std_logic_vector) return int491_t is
  variable rv : int491_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint492_t_to_slv(x : uint492_t) return std_logic_vector is
  variable rv : std_logic_vector(491 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint492_t(x : std_logic_vector) return uint492_t is
  variable rv : uint492_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int492_t_to_slv(x : int492_t) return std_logic_vector is
  variable rv : std_logic_vector(491 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int492_t(x : std_logic_vector) return int492_t is
  variable rv : int492_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint493_t_to_slv(x : uint493_t) return std_logic_vector is
  variable rv : std_logic_vector(492 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint493_t(x : std_logic_vector) return uint493_t is
  variable rv : uint493_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int493_t_to_slv(x : int493_t) return std_logic_vector is
  variable rv : std_logic_vector(492 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int493_t(x : std_logic_vector) return int493_t is
  variable rv : int493_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint494_t_to_slv(x : uint494_t) return std_logic_vector is
  variable rv : std_logic_vector(493 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint494_t(x : std_logic_vector) return uint494_t is
  variable rv : uint494_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int494_t_to_slv(x : int494_t) return std_logic_vector is
  variable rv : std_logic_vector(493 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int494_t(x : std_logic_vector) return int494_t is
  variable rv : int494_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint495_t_to_slv(x : uint495_t) return std_logic_vector is
  variable rv : std_logic_vector(494 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint495_t(x : std_logic_vector) return uint495_t is
  variable rv : uint495_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int495_t_to_slv(x : int495_t) return std_logic_vector is
  variable rv : std_logic_vector(494 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int495_t(x : std_logic_vector) return int495_t is
  variable rv : int495_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint496_t_to_slv(x : uint496_t) return std_logic_vector is
  variable rv : std_logic_vector(495 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint496_t(x : std_logic_vector) return uint496_t is
  variable rv : uint496_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int496_t_to_slv(x : int496_t) return std_logic_vector is
  variable rv : std_logic_vector(495 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int496_t(x : std_logic_vector) return int496_t is
  variable rv : int496_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint497_t_to_slv(x : uint497_t) return std_logic_vector is
  variable rv : std_logic_vector(496 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint497_t(x : std_logic_vector) return uint497_t is
  variable rv : uint497_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int497_t_to_slv(x : int497_t) return std_logic_vector is
  variable rv : std_logic_vector(496 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int497_t(x : std_logic_vector) return int497_t is
  variable rv : int497_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint498_t_to_slv(x : uint498_t) return std_logic_vector is
  variable rv : std_logic_vector(497 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint498_t(x : std_logic_vector) return uint498_t is
  variable rv : uint498_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int498_t_to_slv(x : int498_t) return std_logic_vector is
  variable rv : std_logic_vector(497 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int498_t(x : std_logic_vector) return int498_t is
  variable rv : int498_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint499_t_to_slv(x : uint499_t) return std_logic_vector is
  variable rv : std_logic_vector(498 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint499_t(x : std_logic_vector) return uint499_t is
  variable rv : uint499_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int499_t_to_slv(x : int499_t) return std_logic_vector is
  variable rv : std_logic_vector(498 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int499_t(x : std_logic_vector) return int499_t is
  variable rv : int499_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint500_t_to_slv(x : uint500_t) return std_logic_vector is
  variable rv : std_logic_vector(499 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint500_t(x : std_logic_vector) return uint500_t is
  variable rv : uint500_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int500_t_to_slv(x : int500_t) return std_logic_vector is
  variable rv : std_logic_vector(499 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int500_t(x : std_logic_vector) return int500_t is
  variable rv : int500_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint501_t_to_slv(x : uint501_t) return std_logic_vector is
  variable rv : std_logic_vector(500 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint501_t(x : std_logic_vector) return uint501_t is
  variable rv : uint501_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int501_t_to_slv(x : int501_t) return std_logic_vector is
  variable rv : std_logic_vector(500 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int501_t(x : std_logic_vector) return int501_t is
  variable rv : int501_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint502_t_to_slv(x : uint502_t) return std_logic_vector is
  variable rv : std_logic_vector(501 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint502_t(x : std_logic_vector) return uint502_t is
  variable rv : uint502_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int502_t_to_slv(x : int502_t) return std_logic_vector is
  variable rv : std_logic_vector(501 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int502_t(x : std_logic_vector) return int502_t is
  variable rv : int502_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint503_t_to_slv(x : uint503_t) return std_logic_vector is
  variable rv : std_logic_vector(502 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint503_t(x : std_logic_vector) return uint503_t is
  variable rv : uint503_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int503_t_to_slv(x : int503_t) return std_logic_vector is
  variable rv : std_logic_vector(502 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int503_t(x : std_logic_vector) return int503_t is
  variable rv : int503_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint504_t_to_slv(x : uint504_t) return std_logic_vector is
  variable rv : std_logic_vector(503 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint504_t(x : std_logic_vector) return uint504_t is
  variable rv : uint504_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int504_t_to_slv(x : int504_t) return std_logic_vector is
  variable rv : std_logic_vector(503 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int504_t(x : std_logic_vector) return int504_t is
  variable rv : int504_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint505_t_to_slv(x : uint505_t) return std_logic_vector is
  variable rv : std_logic_vector(504 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint505_t(x : std_logic_vector) return uint505_t is
  variable rv : uint505_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int505_t_to_slv(x : int505_t) return std_logic_vector is
  variable rv : std_logic_vector(504 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int505_t(x : std_logic_vector) return int505_t is
  variable rv : int505_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint506_t_to_slv(x : uint506_t) return std_logic_vector is
  variable rv : std_logic_vector(505 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint506_t(x : std_logic_vector) return uint506_t is
  variable rv : uint506_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int506_t_to_slv(x : int506_t) return std_logic_vector is
  variable rv : std_logic_vector(505 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int506_t(x : std_logic_vector) return int506_t is
  variable rv : int506_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint507_t_to_slv(x : uint507_t) return std_logic_vector is
  variable rv : std_logic_vector(506 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint507_t(x : std_logic_vector) return uint507_t is
  variable rv : uint507_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int507_t_to_slv(x : int507_t) return std_logic_vector is
  variable rv : std_logic_vector(506 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int507_t(x : std_logic_vector) return int507_t is
  variable rv : int507_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint508_t_to_slv(x : uint508_t) return std_logic_vector is
  variable rv : std_logic_vector(507 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint508_t(x : std_logic_vector) return uint508_t is
  variable rv : uint508_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int508_t_to_slv(x : int508_t) return std_logic_vector is
  variable rv : std_logic_vector(507 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int508_t(x : std_logic_vector) return int508_t is
  variable rv : int508_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint509_t_to_slv(x : uint509_t) return std_logic_vector is
  variable rv : std_logic_vector(508 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint509_t(x : std_logic_vector) return uint509_t is
  variable rv : uint509_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int509_t_to_slv(x : int509_t) return std_logic_vector is
  variable rv : std_logic_vector(508 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int509_t(x : std_logic_vector) return int509_t is
  variable rv : int509_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint510_t_to_slv(x : uint510_t) return std_logic_vector is
  variable rv : std_logic_vector(509 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint510_t(x : std_logic_vector) return uint510_t is
  variable rv : uint510_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int510_t_to_slv(x : int510_t) return std_logic_vector is
  variable rv : std_logic_vector(509 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int510_t(x : std_logic_vector) return int510_t is
  variable rv : int510_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint511_t_to_slv(x : uint511_t) return std_logic_vector is
  variable rv : std_logic_vector(510 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint511_t(x : std_logic_vector) return uint511_t is
  variable rv : uint511_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int511_t_to_slv(x : int511_t) return std_logic_vector is
  variable rv : std_logic_vector(510 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int511_t(x : std_logic_vector) return int511_t is
  variable rv : int511_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint512_t_to_slv(x : uint512_t) return std_logic_vector is
  variable rv : std_logic_vector(511 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint512_t(x : std_logic_vector) return uint512_t is
  variable rv : uint512_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int512_t_to_slv(x : int512_t) return std_logic_vector is
  variable rv : std_logic_vector(511 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int512_t(x : std_logic_vector) return int512_t is
  variable rv : int512_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint513_t_to_slv(x : uint513_t) return std_logic_vector is
  variable rv : std_logic_vector(512 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint513_t(x : std_logic_vector) return uint513_t is
  variable rv : uint513_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int513_t_to_slv(x : int513_t) return std_logic_vector is
  variable rv : std_logic_vector(512 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int513_t(x : std_logic_vector) return int513_t is
  variable rv : int513_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint514_t_to_slv(x : uint514_t) return std_logic_vector is
  variable rv : std_logic_vector(513 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint514_t(x : std_logic_vector) return uint514_t is
  variable rv : uint514_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int514_t_to_slv(x : int514_t) return std_logic_vector is
  variable rv : std_logic_vector(513 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int514_t(x : std_logic_vector) return int514_t is
  variable rv : int514_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint515_t_to_slv(x : uint515_t) return std_logic_vector is
  variable rv : std_logic_vector(514 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint515_t(x : std_logic_vector) return uint515_t is
  variable rv : uint515_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int515_t_to_slv(x : int515_t) return std_logic_vector is
  variable rv : std_logic_vector(514 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int515_t(x : std_logic_vector) return int515_t is
  variable rv : int515_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint516_t_to_slv(x : uint516_t) return std_logic_vector is
  variable rv : std_logic_vector(515 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint516_t(x : std_logic_vector) return uint516_t is
  variable rv : uint516_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int516_t_to_slv(x : int516_t) return std_logic_vector is
  variable rv : std_logic_vector(515 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int516_t(x : std_logic_vector) return int516_t is
  variable rv : int516_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint517_t_to_slv(x : uint517_t) return std_logic_vector is
  variable rv : std_logic_vector(516 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint517_t(x : std_logic_vector) return uint517_t is
  variable rv : uint517_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int517_t_to_slv(x : int517_t) return std_logic_vector is
  variable rv : std_logic_vector(516 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int517_t(x : std_logic_vector) return int517_t is
  variable rv : int517_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint518_t_to_slv(x : uint518_t) return std_logic_vector is
  variable rv : std_logic_vector(517 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint518_t(x : std_logic_vector) return uint518_t is
  variable rv : uint518_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int518_t_to_slv(x : int518_t) return std_logic_vector is
  variable rv : std_logic_vector(517 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int518_t(x : std_logic_vector) return int518_t is
  variable rv : int518_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint519_t_to_slv(x : uint519_t) return std_logic_vector is
  variable rv : std_logic_vector(518 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint519_t(x : std_logic_vector) return uint519_t is
  variable rv : uint519_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int519_t_to_slv(x : int519_t) return std_logic_vector is
  variable rv : std_logic_vector(518 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int519_t(x : std_logic_vector) return int519_t is
  variable rv : int519_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint520_t_to_slv(x : uint520_t) return std_logic_vector is
  variable rv : std_logic_vector(519 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint520_t(x : std_logic_vector) return uint520_t is
  variable rv : uint520_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int520_t_to_slv(x : int520_t) return std_logic_vector is
  variable rv : std_logic_vector(519 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int520_t(x : std_logic_vector) return int520_t is
  variable rv : int520_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint521_t_to_slv(x : uint521_t) return std_logic_vector is
  variable rv : std_logic_vector(520 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint521_t(x : std_logic_vector) return uint521_t is
  variable rv : uint521_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int521_t_to_slv(x : int521_t) return std_logic_vector is
  variable rv : std_logic_vector(520 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int521_t(x : std_logic_vector) return int521_t is
  variable rv : int521_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint522_t_to_slv(x : uint522_t) return std_logic_vector is
  variable rv : std_logic_vector(521 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint522_t(x : std_logic_vector) return uint522_t is
  variable rv : uint522_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int522_t_to_slv(x : int522_t) return std_logic_vector is
  variable rv : std_logic_vector(521 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int522_t(x : std_logic_vector) return int522_t is
  variable rv : int522_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint523_t_to_slv(x : uint523_t) return std_logic_vector is
  variable rv : std_logic_vector(522 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint523_t(x : std_logic_vector) return uint523_t is
  variable rv : uint523_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int523_t_to_slv(x : int523_t) return std_logic_vector is
  variable rv : std_logic_vector(522 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int523_t(x : std_logic_vector) return int523_t is
  variable rv : int523_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint524_t_to_slv(x : uint524_t) return std_logic_vector is
  variable rv : std_logic_vector(523 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint524_t(x : std_logic_vector) return uint524_t is
  variable rv : uint524_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int524_t_to_slv(x : int524_t) return std_logic_vector is
  variable rv : std_logic_vector(523 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int524_t(x : std_logic_vector) return int524_t is
  variable rv : int524_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint525_t_to_slv(x : uint525_t) return std_logic_vector is
  variable rv : std_logic_vector(524 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint525_t(x : std_logic_vector) return uint525_t is
  variable rv : uint525_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int525_t_to_slv(x : int525_t) return std_logic_vector is
  variable rv : std_logic_vector(524 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int525_t(x : std_logic_vector) return int525_t is
  variable rv : int525_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint526_t_to_slv(x : uint526_t) return std_logic_vector is
  variable rv : std_logic_vector(525 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint526_t(x : std_logic_vector) return uint526_t is
  variable rv : uint526_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int526_t_to_slv(x : int526_t) return std_logic_vector is
  variable rv : std_logic_vector(525 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int526_t(x : std_logic_vector) return int526_t is
  variable rv : int526_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint527_t_to_slv(x : uint527_t) return std_logic_vector is
  variable rv : std_logic_vector(526 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint527_t(x : std_logic_vector) return uint527_t is
  variable rv : uint527_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int527_t_to_slv(x : int527_t) return std_logic_vector is
  variable rv : std_logic_vector(526 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int527_t(x : std_logic_vector) return int527_t is
  variable rv : int527_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint528_t_to_slv(x : uint528_t) return std_logic_vector is
  variable rv : std_logic_vector(527 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint528_t(x : std_logic_vector) return uint528_t is
  variable rv : uint528_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int528_t_to_slv(x : int528_t) return std_logic_vector is
  variable rv : std_logic_vector(527 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int528_t(x : std_logic_vector) return int528_t is
  variable rv : int528_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint529_t_to_slv(x : uint529_t) return std_logic_vector is
  variable rv : std_logic_vector(528 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint529_t(x : std_logic_vector) return uint529_t is
  variable rv : uint529_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int529_t_to_slv(x : int529_t) return std_logic_vector is
  variable rv : std_logic_vector(528 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int529_t(x : std_logic_vector) return int529_t is
  variable rv : int529_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint530_t_to_slv(x : uint530_t) return std_logic_vector is
  variable rv : std_logic_vector(529 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint530_t(x : std_logic_vector) return uint530_t is
  variable rv : uint530_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int530_t_to_slv(x : int530_t) return std_logic_vector is
  variable rv : std_logic_vector(529 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int530_t(x : std_logic_vector) return int530_t is
  variable rv : int530_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint531_t_to_slv(x : uint531_t) return std_logic_vector is
  variable rv : std_logic_vector(530 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint531_t(x : std_logic_vector) return uint531_t is
  variable rv : uint531_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int531_t_to_slv(x : int531_t) return std_logic_vector is
  variable rv : std_logic_vector(530 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int531_t(x : std_logic_vector) return int531_t is
  variable rv : int531_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint532_t_to_slv(x : uint532_t) return std_logic_vector is
  variable rv : std_logic_vector(531 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint532_t(x : std_logic_vector) return uint532_t is
  variable rv : uint532_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int532_t_to_slv(x : int532_t) return std_logic_vector is
  variable rv : std_logic_vector(531 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int532_t(x : std_logic_vector) return int532_t is
  variable rv : int532_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint533_t_to_slv(x : uint533_t) return std_logic_vector is
  variable rv : std_logic_vector(532 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint533_t(x : std_logic_vector) return uint533_t is
  variable rv : uint533_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int533_t_to_slv(x : int533_t) return std_logic_vector is
  variable rv : std_logic_vector(532 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int533_t(x : std_logic_vector) return int533_t is
  variable rv : int533_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint534_t_to_slv(x : uint534_t) return std_logic_vector is
  variable rv : std_logic_vector(533 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint534_t(x : std_logic_vector) return uint534_t is
  variable rv : uint534_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int534_t_to_slv(x : int534_t) return std_logic_vector is
  variable rv : std_logic_vector(533 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int534_t(x : std_logic_vector) return int534_t is
  variable rv : int534_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint535_t_to_slv(x : uint535_t) return std_logic_vector is
  variable rv : std_logic_vector(534 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint535_t(x : std_logic_vector) return uint535_t is
  variable rv : uint535_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int535_t_to_slv(x : int535_t) return std_logic_vector is
  variable rv : std_logic_vector(534 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int535_t(x : std_logic_vector) return int535_t is
  variable rv : int535_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint536_t_to_slv(x : uint536_t) return std_logic_vector is
  variable rv : std_logic_vector(535 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint536_t(x : std_logic_vector) return uint536_t is
  variable rv : uint536_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int536_t_to_slv(x : int536_t) return std_logic_vector is
  variable rv : std_logic_vector(535 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int536_t(x : std_logic_vector) return int536_t is
  variable rv : int536_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint537_t_to_slv(x : uint537_t) return std_logic_vector is
  variable rv : std_logic_vector(536 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint537_t(x : std_logic_vector) return uint537_t is
  variable rv : uint537_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int537_t_to_slv(x : int537_t) return std_logic_vector is
  variable rv : std_logic_vector(536 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int537_t(x : std_logic_vector) return int537_t is
  variable rv : int537_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint538_t_to_slv(x : uint538_t) return std_logic_vector is
  variable rv : std_logic_vector(537 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint538_t(x : std_logic_vector) return uint538_t is
  variable rv : uint538_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int538_t_to_slv(x : int538_t) return std_logic_vector is
  variable rv : std_logic_vector(537 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int538_t(x : std_logic_vector) return int538_t is
  variable rv : int538_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint539_t_to_slv(x : uint539_t) return std_logic_vector is
  variable rv : std_logic_vector(538 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint539_t(x : std_logic_vector) return uint539_t is
  variable rv : uint539_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int539_t_to_slv(x : int539_t) return std_logic_vector is
  variable rv : std_logic_vector(538 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int539_t(x : std_logic_vector) return int539_t is
  variable rv : int539_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint540_t_to_slv(x : uint540_t) return std_logic_vector is
  variable rv : std_logic_vector(539 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint540_t(x : std_logic_vector) return uint540_t is
  variable rv : uint540_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int540_t_to_slv(x : int540_t) return std_logic_vector is
  variable rv : std_logic_vector(539 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int540_t(x : std_logic_vector) return int540_t is
  variable rv : int540_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint541_t_to_slv(x : uint541_t) return std_logic_vector is
  variable rv : std_logic_vector(540 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint541_t(x : std_logic_vector) return uint541_t is
  variable rv : uint541_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int541_t_to_slv(x : int541_t) return std_logic_vector is
  variable rv : std_logic_vector(540 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int541_t(x : std_logic_vector) return int541_t is
  variable rv : int541_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint542_t_to_slv(x : uint542_t) return std_logic_vector is
  variable rv : std_logic_vector(541 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint542_t(x : std_logic_vector) return uint542_t is
  variable rv : uint542_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int542_t_to_slv(x : int542_t) return std_logic_vector is
  variable rv : std_logic_vector(541 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int542_t(x : std_logic_vector) return int542_t is
  variable rv : int542_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint543_t_to_slv(x : uint543_t) return std_logic_vector is
  variable rv : std_logic_vector(542 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint543_t(x : std_logic_vector) return uint543_t is
  variable rv : uint543_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int543_t_to_slv(x : int543_t) return std_logic_vector is
  variable rv : std_logic_vector(542 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int543_t(x : std_logic_vector) return int543_t is
  variable rv : int543_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint544_t_to_slv(x : uint544_t) return std_logic_vector is
  variable rv : std_logic_vector(543 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint544_t(x : std_logic_vector) return uint544_t is
  variable rv : uint544_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int544_t_to_slv(x : int544_t) return std_logic_vector is
  variable rv : std_logic_vector(543 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int544_t(x : std_logic_vector) return int544_t is
  variable rv : int544_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint545_t_to_slv(x : uint545_t) return std_logic_vector is
  variable rv : std_logic_vector(544 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint545_t(x : std_logic_vector) return uint545_t is
  variable rv : uint545_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int545_t_to_slv(x : int545_t) return std_logic_vector is
  variable rv : std_logic_vector(544 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int545_t(x : std_logic_vector) return int545_t is
  variable rv : int545_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint546_t_to_slv(x : uint546_t) return std_logic_vector is
  variable rv : std_logic_vector(545 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint546_t(x : std_logic_vector) return uint546_t is
  variable rv : uint546_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int546_t_to_slv(x : int546_t) return std_logic_vector is
  variable rv : std_logic_vector(545 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int546_t(x : std_logic_vector) return int546_t is
  variable rv : int546_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint547_t_to_slv(x : uint547_t) return std_logic_vector is
  variable rv : std_logic_vector(546 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint547_t(x : std_logic_vector) return uint547_t is
  variable rv : uint547_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int547_t_to_slv(x : int547_t) return std_logic_vector is
  variable rv : std_logic_vector(546 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int547_t(x : std_logic_vector) return int547_t is
  variable rv : int547_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint548_t_to_slv(x : uint548_t) return std_logic_vector is
  variable rv : std_logic_vector(547 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint548_t(x : std_logic_vector) return uint548_t is
  variable rv : uint548_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int548_t_to_slv(x : int548_t) return std_logic_vector is
  variable rv : std_logic_vector(547 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int548_t(x : std_logic_vector) return int548_t is
  variable rv : int548_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint549_t_to_slv(x : uint549_t) return std_logic_vector is
  variable rv : std_logic_vector(548 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint549_t(x : std_logic_vector) return uint549_t is
  variable rv : uint549_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int549_t_to_slv(x : int549_t) return std_logic_vector is
  variable rv : std_logic_vector(548 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int549_t(x : std_logic_vector) return int549_t is
  variable rv : int549_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint550_t_to_slv(x : uint550_t) return std_logic_vector is
  variable rv : std_logic_vector(549 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint550_t(x : std_logic_vector) return uint550_t is
  variable rv : uint550_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int550_t_to_slv(x : int550_t) return std_logic_vector is
  variable rv : std_logic_vector(549 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int550_t(x : std_logic_vector) return int550_t is
  variable rv : int550_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint551_t_to_slv(x : uint551_t) return std_logic_vector is
  variable rv : std_logic_vector(550 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint551_t(x : std_logic_vector) return uint551_t is
  variable rv : uint551_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int551_t_to_slv(x : int551_t) return std_logic_vector is
  variable rv : std_logic_vector(550 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int551_t(x : std_logic_vector) return int551_t is
  variable rv : int551_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint552_t_to_slv(x : uint552_t) return std_logic_vector is
  variable rv : std_logic_vector(551 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint552_t(x : std_logic_vector) return uint552_t is
  variable rv : uint552_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int552_t_to_slv(x : int552_t) return std_logic_vector is
  variable rv : std_logic_vector(551 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int552_t(x : std_logic_vector) return int552_t is
  variable rv : int552_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint553_t_to_slv(x : uint553_t) return std_logic_vector is
  variable rv : std_logic_vector(552 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint553_t(x : std_logic_vector) return uint553_t is
  variable rv : uint553_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int553_t_to_slv(x : int553_t) return std_logic_vector is
  variable rv : std_logic_vector(552 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int553_t(x : std_logic_vector) return int553_t is
  variable rv : int553_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint554_t_to_slv(x : uint554_t) return std_logic_vector is
  variable rv : std_logic_vector(553 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint554_t(x : std_logic_vector) return uint554_t is
  variable rv : uint554_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int554_t_to_slv(x : int554_t) return std_logic_vector is
  variable rv : std_logic_vector(553 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int554_t(x : std_logic_vector) return int554_t is
  variable rv : int554_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint555_t_to_slv(x : uint555_t) return std_logic_vector is
  variable rv : std_logic_vector(554 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint555_t(x : std_logic_vector) return uint555_t is
  variable rv : uint555_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int555_t_to_slv(x : int555_t) return std_logic_vector is
  variable rv : std_logic_vector(554 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int555_t(x : std_logic_vector) return int555_t is
  variable rv : int555_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint556_t_to_slv(x : uint556_t) return std_logic_vector is
  variable rv : std_logic_vector(555 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint556_t(x : std_logic_vector) return uint556_t is
  variable rv : uint556_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int556_t_to_slv(x : int556_t) return std_logic_vector is
  variable rv : std_logic_vector(555 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int556_t(x : std_logic_vector) return int556_t is
  variable rv : int556_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint557_t_to_slv(x : uint557_t) return std_logic_vector is
  variable rv : std_logic_vector(556 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint557_t(x : std_logic_vector) return uint557_t is
  variable rv : uint557_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int557_t_to_slv(x : int557_t) return std_logic_vector is
  variable rv : std_logic_vector(556 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int557_t(x : std_logic_vector) return int557_t is
  variable rv : int557_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint558_t_to_slv(x : uint558_t) return std_logic_vector is
  variable rv : std_logic_vector(557 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint558_t(x : std_logic_vector) return uint558_t is
  variable rv : uint558_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int558_t_to_slv(x : int558_t) return std_logic_vector is
  variable rv : std_logic_vector(557 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int558_t(x : std_logic_vector) return int558_t is
  variable rv : int558_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint559_t_to_slv(x : uint559_t) return std_logic_vector is
  variable rv : std_logic_vector(558 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint559_t(x : std_logic_vector) return uint559_t is
  variable rv : uint559_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int559_t_to_slv(x : int559_t) return std_logic_vector is
  variable rv : std_logic_vector(558 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int559_t(x : std_logic_vector) return int559_t is
  variable rv : int559_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint560_t_to_slv(x : uint560_t) return std_logic_vector is
  variable rv : std_logic_vector(559 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint560_t(x : std_logic_vector) return uint560_t is
  variable rv : uint560_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int560_t_to_slv(x : int560_t) return std_logic_vector is
  variable rv : std_logic_vector(559 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int560_t(x : std_logic_vector) return int560_t is
  variable rv : int560_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint561_t_to_slv(x : uint561_t) return std_logic_vector is
  variable rv : std_logic_vector(560 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint561_t(x : std_logic_vector) return uint561_t is
  variable rv : uint561_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int561_t_to_slv(x : int561_t) return std_logic_vector is
  variable rv : std_logic_vector(560 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int561_t(x : std_logic_vector) return int561_t is
  variable rv : int561_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint562_t_to_slv(x : uint562_t) return std_logic_vector is
  variable rv : std_logic_vector(561 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint562_t(x : std_logic_vector) return uint562_t is
  variable rv : uint562_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int562_t_to_slv(x : int562_t) return std_logic_vector is
  variable rv : std_logic_vector(561 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int562_t(x : std_logic_vector) return int562_t is
  variable rv : int562_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint563_t_to_slv(x : uint563_t) return std_logic_vector is
  variable rv : std_logic_vector(562 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint563_t(x : std_logic_vector) return uint563_t is
  variable rv : uint563_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int563_t_to_slv(x : int563_t) return std_logic_vector is
  variable rv : std_logic_vector(562 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int563_t(x : std_logic_vector) return int563_t is
  variable rv : int563_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint564_t_to_slv(x : uint564_t) return std_logic_vector is
  variable rv : std_logic_vector(563 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint564_t(x : std_logic_vector) return uint564_t is
  variable rv : uint564_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int564_t_to_slv(x : int564_t) return std_logic_vector is
  variable rv : std_logic_vector(563 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int564_t(x : std_logic_vector) return int564_t is
  variable rv : int564_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint565_t_to_slv(x : uint565_t) return std_logic_vector is
  variable rv : std_logic_vector(564 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint565_t(x : std_logic_vector) return uint565_t is
  variable rv : uint565_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int565_t_to_slv(x : int565_t) return std_logic_vector is
  variable rv : std_logic_vector(564 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int565_t(x : std_logic_vector) return int565_t is
  variable rv : int565_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint566_t_to_slv(x : uint566_t) return std_logic_vector is
  variable rv : std_logic_vector(565 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint566_t(x : std_logic_vector) return uint566_t is
  variable rv : uint566_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int566_t_to_slv(x : int566_t) return std_logic_vector is
  variable rv : std_logic_vector(565 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int566_t(x : std_logic_vector) return int566_t is
  variable rv : int566_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint567_t_to_slv(x : uint567_t) return std_logic_vector is
  variable rv : std_logic_vector(566 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint567_t(x : std_logic_vector) return uint567_t is
  variable rv : uint567_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int567_t_to_slv(x : int567_t) return std_logic_vector is
  variable rv : std_logic_vector(566 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int567_t(x : std_logic_vector) return int567_t is
  variable rv : int567_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint568_t_to_slv(x : uint568_t) return std_logic_vector is
  variable rv : std_logic_vector(567 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint568_t(x : std_logic_vector) return uint568_t is
  variable rv : uint568_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int568_t_to_slv(x : int568_t) return std_logic_vector is
  variable rv : std_logic_vector(567 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int568_t(x : std_logic_vector) return int568_t is
  variable rv : int568_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint569_t_to_slv(x : uint569_t) return std_logic_vector is
  variable rv : std_logic_vector(568 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint569_t(x : std_logic_vector) return uint569_t is
  variable rv : uint569_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int569_t_to_slv(x : int569_t) return std_logic_vector is
  variable rv : std_logic_vector(568 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int569_t(x : std_logic_vector) return int569_t is
  variable rv : int569_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint570_t_to_slv(x : uint570_t) return std_logic_vector is
  variable rv : std_logic_vector(569 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint570_t(x : std_logic_vector) return uint570_t is
  variable rv : uint570_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int570_t_to_slv(x : int570_t) return std_logic_vector is
  variable rv : std_logic_vector(569 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int570_t(x : std_logic_vector) return int570_t is
  variable rv : int570_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint571_t_to_slv(x : uint571_t) return std_logic_vector is
  variable rv : std_logic_vector(570 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint571_t(x : std_logic_vector) return uint571_t is
  variable rv : uint571_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int571_t_to_slv(x : int571_t) return std_logic_vector is
  variable rv : std_logic_vector(570 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int571_t(x : std_logic_vector) return int571_t is
  variable rv : int571_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint572_t_to_slv(x : uint572_t) return std_logic_vector is
  variable rv : std_logic_vector(571 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint572_t(x : std_logic_vector) return uint572_t is
  variable rv : uint572_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int572_t_to_slv(x : int572_t) return std_logic_vector is
  variable rv : std_logic_vector(571 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int572_t(x : std_logic_vector) return int572_t is
  variable rv : int572_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint573_t_to_slv(x : uint573_t) return std_logic_vector is
  variable rv : std_logic_vector(572 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint573_t(x : std_logic_vector) return uint573_t is
  variable rv : uint573_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int573_t_to_slv(x : int573_t) return std_logic_vector is
  variable rv : std_logic_vector(572 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int573_t(x : std_logic_vector) return int573_t is
  variable rv : int573_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint574_t_to_slv(x : uint574_t) return std_logic_vector is
  variable rv : std_logic_vector(573 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint574_t(x : std_logic_vector) return uint574_t is
  variable rv : uint574_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int574_t_to_slv(x : int574_t) return std_logic_vector is
  variable rv : std_logic_vector(573 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int574_t(x : std_logic_vector) return int574_t is
  variable rv : int574_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint575_t_to_slv(x : uint575_t) return std_logic_vector is
  variable rv : std_logic_vector(574 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint575_t(x : std_logic_vector) return uint575_t is
  variable rv : uint575_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int575_t_to_slv(x : int575_t) return std_logic_vector is
  variable rv : std_logic_vector(574 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int575_t(x : std_logic_vector) return int575_t is
  variable rv : int575_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint576_t_to_slv(x : uint576_t) return std_logic_vector is
  variable rv : std_logic_vector(575 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint576_t(x : std_logic_vector) return uint576_t is
  variable rv : uint576_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int576_t_to_slv(x : int576_t) return std_logic_vector is
  variable rv : std_logic_vector(575 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int576_t(x : std_logic_vector) return int576_t is
  variable rv : int576_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint577_t_to_slv(x : uint577_t) return std_logic_vector is
  variable rv : std_logic_vector(576 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint577_t(x : std_logic_vector) return uint577_t is
  variable rv : uint577_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int577_t_to_slv(x : int577_t) return std_logic_vector is
  variable rv : std_logic_vector(576 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int577_t(x : std_logic_vector) return int577_t is
  variable rv : int577_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint578_t_to_slv(x : uint578_t) return std_logic_vector is
  variable rv : std_logic_vector(577 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint578_t(x : std_logic_vector) return uint578_t is
  variable rv : uint578_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int578_t_to_slv(x : int578_t) return std_logic_vector is
  variable rv : std_logic_vector(577 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int578_t(x : std_logic_vector) return int578_t is
  variable rv : int578_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint579_t_to_slv(x : uint579_t) return std_logic_vector is
  variable rv : std_logic_vector(578 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint579_t(x : std_logic_vector) return uint579_t is
  variable rv : uint579_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int579_t_to_slv(x : int579_t) return std_logic_vector is
  variable rv : std_logic_vector(578 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int579_t(x : std_logic_vector) return int579_t is
  variable rv : int579_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint580_t_to_slv(x : uint580_t) return std_logic_vector is
  variable rv : std_logic_vector(579 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint580_t(x : std_logic_vector) return uint580_t is
  variable rv : uint580_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int580_t_to_slv(x : int580_t) return std_logic_vector is
  variable rv : std_logic_vector(579 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int580_t(x : std_logic_vector) return int580_t is
  variable rv : int580_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint581_t_to_slv(x : uint581_t) return std_logic_vector is
  variable rv : std_logic_vector(580 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint581_t(x : std_logic_vector) return uint581_t is
  variable rv : uint581_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int581_t_to_slv(x : int581_t) return std_logic_vector is
  variable rv : std_logic_vector(580 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int581_t(x : std_logic_vector) return int581_t is
  variable rv : int581_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint582_t_to_slv(x : uint582_t) return std_logic_vector is
  variable rv : std_logic_vector(581 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint582_t(x : std_logic_vector) return uint582_t is
  variable rv : uint582_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int582_t_to_slv(x : int582_t) return std_logic_vector is
  variable rv : std_logic_vector(581 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int582_t(x : std_logic_vector) return int582_t is
  variable rv : int582_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint583_t_to_slv(x : uint583_t) return std_logic_vector is
  variable rv : std_logic_vector(582 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint583_t(x : std_logic_vector) return uint583_t is
  variable rv : uint583_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int583_t_to_slv(x : int583_t) return std_logic_vector is
  variable rv : std_logic_vector(582 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int583_t(x : std_logic_vector) return int583_t is
  variable rv : int583_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint584_t_to_slv(x : uint584_t) return std_logic_vector is
  variable rv : std_logic_vector(583 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint584_t(x : std_logic_vector) return uint584_t is
  variable rv : uint584_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int584_t_to_slv(x : int584_t) return std_logic_vector is
  variable rv : std_logic_vector(583 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int584_t(x : std_logic_vector) return int584_t is
  variable rv : int584_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint585_t_to_slv(x : uint585_t) return std_logic_vector is
  variable rv : std_logic_vector(584 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint585_t(x : std_logic_vector) return uint585_t is
  variable rv : uint585_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int585_t_to_slv(x : int585_t) return std_logic_vector is
  variable rv : std_logic_vector(584 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int585_t(x : std_logic_vector) return int585_t is
  variable rv : int585_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint586_t_to_slv(x : uint586_t) return std_logic_vector is
  variable rv : std_logic_vector(585 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint586_t(x : std_logic_vector) return uint586_t is
  variable rv : uint586_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int586_t_to_slv(x : int586_t) return std_logic_vector is
  variable rv : std_logic_vector(585 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int586_t(x : std_logic_vector) return int586_t is
  variable rv : int586_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint587_t_to_slv(x : uint587_t) return std_logic_vector is
  variable rv : std_logic_vector(586 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint587_t(x : std_logic_vector) return uint587_t is
  variable rv : uint587_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int587_t_to_slv(x : int587_t) return std_logic_vector is
  variable rv : std_logic_vector(586 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int587_t(x : std_logic_vector) return int587_t is
  variable rv : int587_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint588_t_to_slv(x : uint588_t) return std_logic_vector is
  variable rv : std_logic_vector(587 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint588_t(x : std_logic_vector) return uint588_t is
  variable rv : uint588_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int588_t_to_slv(x : int588_t) return std_logic_vector is
  variable rv : std_logic_vector(587 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int588_t(x : std_logic_vector) return int588_t is
  variable rv : int588_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint589_t_to_slv(x : uint589_t) return std_logic_vector is
  variable rv : std_logic_vector(588 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint589_t(x : std_logic_vector) return uint589_t is
  variable rv : uint589_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int589_t_to_slv(x : int589_t) return std_logic_vector is
  variable rv : std_logic_vector(588 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int589_t(x : std_logic_vector) return int589_t is
  variable rv : int589_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint590_t_to_slv(x : uint590_t) return std_logic_vector is
  variable rv : std_logic_vector(589 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint590_t(x : std_logic_vector) return uint590_t is
  variable rv : uint590_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int590_t_to_slv(x : int590_t) return std_logic_vector is
  variable rv : std_logic_vector(589 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int590_t(x : std_logic_vector) return int590_t is
  variable rv : int590_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint591_t_to_slv(x : uint591_t) return std_logic_vector is
  variable rv : std_logic_vector(590 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint591_t(x : std_logic_vector) return uint591_t is
  variable rv : uint591_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int591_t_to_slv(x : int591_t) return std_logic_vector is
  variable rv : std_logic_vector(590 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int591_t(x : std_logic_vector) return int591_t is
  variable rv : int591_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint592_t_to_slv(x : uint592_t) return std_logic_vector is
  variable rv : std_logic_vector(591 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint592_t(x : std_logic_vector) return uint592_t is
  variable rv : uint592_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int592_t_to_slv(x : int592_t) return std_logic_vector is
  variable rv : std_logic_vector(591 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int592_t(x : std_logic_vector) return int592_t is
  variable rv : int592_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint593_t_to_slv(x : uint593_t) return std_logic_vector is
  variable rv : std_logic_vector(592 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint593_t(x : std_logic_vector) return uint593_t is
  variable rv : uint593_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int593_t_to_slv(x : int593_t) return std_logic_vector is
  variable rv : std_logic_vector(592 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int593_t(x : std_logic_vector) return int593_t is
  variable rv : int593_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint594_t_to_slv(x : uint594_t) return std_logic_vector is
  variable rv : std_logic_vector(593 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint594_t(x : std_logic_vector) return uint594_t is
  variable rv : uint594_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int594_t_to_slv(x : int594_t) return std_logic_vector is
  variable rv : std_logic_vector(593 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int594_t(x : std_logic_vector) return int594_t is
  variable rv : int594_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint595_t_to_slv(x : uint595_t) return std_logic_vector is
  variable rv : std_logic_vector(594 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint595_t(x : std_logic_vector) return uint595_t is
  variable rv : uint595_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int595_t_to_slv(x : int595_t) return std_logic_vector is
  variable rv : std_logic_vector(594 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int595_t(x : std_logic_vector) return int595_t is
  variable rv : int595_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint596_t_to_slv(x : uint596_t) return std_logic_vector is
  variable rv : std_logic_vector(595 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint596_t(x : std_logic_vector) return uint596_t is
  variable rv : uint596_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int596_t_to_slv(x : int596_t) return std_logic_vector is
  variable rv : std_logic_vector(595 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int596_t(x : std_logic_vector) return int596_t is
  variable rv : int596_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint597_t_to_slv(x : uint597_t) return std_logic_vector is
  variable rv : std_logic_vector(596 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint597_t(x : std_logic_vector) return uint597_t is
  variable rv : uint597_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int597_t_to_slv(x : int597_t) return std_logic_vector is
  variable rv : std_logic_vector(596 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int597_t(x : std_logic_vector) return int597_t is
  variable rv : int597_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint598_t_to_slv(x : uint598_t) return std_logic_vector is
  variable rv : std_logic_vector(597 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint598_t(x : std_logic_vector) return uint598_t is
  variable rv : uint598_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int598_t_to_slv(x : int598_t) return std_logic_vector is
  variable rv : std_logic_vector(597 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int598_t(x : std_logic_vector) return int598_t is
  variable rv : int598_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint599_t_to_slv(x : uint599_t) return std_logic_vector is
  variable rv : std_logic_vector(598 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint599_t(x : std_logic_vector) return uint599_t is
  variable rv : uint599_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int599_t_to_slv(x : int599_t) return std_logic_vector is
  variable rv : std_logic_vector(598 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int599_t(x : std_logic_vector) return int599_t is
  variable rv : int599_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint600_t_to_slv(x : uint600_t) return std_logic_vector is
  variable rv : std_logic_vector(599 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint600_t(x : std_logic_vector) return uint600_t is
  variable rv : uint600_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int600_t_to_slv(x : int600_t) return std_logic_vector is
  variable rv : std_logic_vector(599 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int600_t(x : std_logic_vector) return int600_t is
  variable rv : int600_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint601_t_to_slv(x : uint601_t) return std_logic_vector is
  variable rv : std_logic_vector(600 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint601_t(x : std_logic_vector) return uint601_t is
  variable rv : uint601_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int601_t_to_slv(x : int601_t) return std_logic_vector is
  variable rv : std_logic_vector(600 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int601_t(x : std_logic_vector) return int601_t is
  variable rv : int601_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint602_t_to_slv(x : uint602_t) return std_logic_vector is
  variable rv : std_logic_vector(601 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint602_t(x : std_logic_vector) return uint602_t is
  variable rv : uint602_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int602_t_to_slv(x : int602_t) return std_logic_vector is
  variable rv : std_logic_vector(601 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int602_t(x : std_logic_vector) return int602_t is
  variable rv : int602_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint603_t_to_slv(x : uint603_t) return std_logic_vector is
  variable rv : std_logic_vector(602 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint603_t(x : std_logic_vector) return uint603_t is
  variable rv : uint603_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int603_t_to_slv(x : int603_t) return std_logic_vector is
  variable rv : std_logic_vector(602 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int603_t(x : std_logic_vector) return int603_t is
  variable rv : int603_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint604_t_to_slv(x : uint604_t) return std_logic_vector is
  variable rv : std_logic_vector(603 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint604_t(x : std_logic_vector) return uint604_t is
  variable rv : uint604_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int604_t_to_slv(x : int604_t) return std_logic_vector is
  variable rv : std_logic_vector(603 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int604_t(x : std_logic_vector) return int604_t is
  variable rv : int604_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint605_t_to_slv(x : uint605_t) return std_logic_vector is
  variable rv : std_logic_vector(604 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint605_t(x : std_logic_vector) return uint605_t is
  variable rv : uint605_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int605_t_to_slv(x : int605_t) return std_logic_vector is
  variable rv : std_logic_vector(604 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int605_t(x : std_logic_vector) return int605_t is
  variable rv : int605_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint606_t_to_slv(x : uint606_t) return std_logic_vector is
  variable rv : std_logic_vector(605 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint606_t(x : std_logic_vector) return uint606_t is
  variable rv : uint606_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int606_t_to_slv(x : int606_t) return std_logic_vector is
  variable rv : std_logic_vector(605 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int606_t(x : std_logic_vector) return int606_t is
  variable rv : int606_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint607_t_to_slv(x : uint607_t) return std_logic_vector is
  variable rv : std_logic_vector(606 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint607_t(x : std_logic_vector) return uint607_t is
  variable rv : uint607_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int607_t_to_slv(x : int607_t) return std_logic_vector is
  variable rv : std_logic_vector(606 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int607_t(x : std_logic_vector) return int607_t is
  variable rv : int607_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint608_t_to_slv(x : uint608_t) return std_logic_vector is
  variable rv : std_logic_vector(607 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint608_t(x : std_logic_vector) return uint608_t is
  variable rv : uint608_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int608_t_to_slv(x : int608_t) return std_logic_vector is
  variable rv : std_logic_vector(607 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int608_t(x : std_logic_vector) return int608_t is
  variable rv : int608_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint609_t_to_slv(x : uint609_t) return std_logic_vector is
  variable rv : std_logic_vector(608 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint609_t(x : std_logic_vector) return uint609_t is
  variable rv : uint609_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int609_t_to_slv(x : int609_t) return std_logic_vector is
  variable rv : std_logic_vector(608 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int609_t(x : std_logic_vector) return int609_t is
  variable rv : int609_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint610_t_to_slv(x : uint610_t) return std_logic_vector is
  variable rv : std_logic_vector(609 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint610_t(x : std_logic_vector) return uint610_t is
  variable rv : uint610_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int610_t_to_slv(x : int610_t) return std_logic_vector is
  variable rv : std_logic_vector(609 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int610_t(x : std_logic_vector) return int610_t is
  variable rv : int610_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint611_t_to_slv(x : uint611_t) return std_logic_vector is
  variable rv : std_logic_vector(610 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint611_t(x : std_logic_vector) return uint611_t is
  variable rv : uint611_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int611_t_to_slv(x : int611_t) return std_logic_vector is
  variable rv : std_logic_vector(610 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int611_t(x : std_logic_vector) return int611_t is
  variable rv : int611_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint612_t_to_slv(x : uint612_t) return std_logic_vector is
  variable rv : std_logic_vector(611 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint612_t(x : std_logic_vector) return uint612_t is
  variable rv : uint612_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int612_t_to_slv(x : int612_t) return std_logic_vector is
  variable rv : std_logic_vector(611 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int612_t(x : std_logic_vector) return int612_t is
  variable rv : int612_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint613_t_to_slv(x : uint613_t) return std_logic_vector is
  variable rv : std_logic_vector(612 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint613_t(x : std_logic_vector) return uint613_t is
  variable rv : uint613_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int613_t_to_slv(x : int613_t) return std_logic_vector is
  variable rv : std_logic_vector(612 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int613_t(x : std_logic_vector) return int613_t is
  variable rv : int613_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint614_t_to_slv(x : uint614_t) return std_logic_vector is
  variable rv : std_logic_vector(613 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint614_t(x : std_logic_vector) return uint614_t is
  variable rv : uint614_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int614_t_to_slv(x : int614_t) return std_logic_vector is
  variable rv : std_logic_vector(613 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int614_t(x : std_logic_vector) return int614_t is
  variable rv : int614_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint615_t_to_slv(x : uint615_t) return std_logic_vector is
  variable rv : std_logic_vector(614 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint615_t(x : std_logic_vector) return uint615_t is
  variable rv : uint615_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int615_t_to_slv(x : int615_t) return std_logic_vector is
  variable rv : std_logic_vector(614 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int615_t(x : std_logic_vector) return int615_t is
  variable rv : int615_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint616_t_to_slv(x : uint616_t) return std_logic_vector is
  variable rv : std_logic_vector(615 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint616_t(x : std_logic_vector) return uint616_t is
  variable rv : uint616_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int616_t_to_slv(x : int616_t) return std_logic_vector is
  variable rv : std_logic_vector(615 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int616_t(x : std_logic_vector) return int616_t is
  variable rv : int616_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint617_t_to_slv(x : uint617_t) return std_logic_vector is
  variable rv : std_logic_vector(616 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint617_t(x : std_logic_vector) return uint617_t is
  variable rv : uint617_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int617_t_to_slv(x : int617_t) return std_logic_vector is
  variable rv : std_logic_vector(616 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int617_t(x : std_logic_vector) return int617_t is
  variable rv : int617_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint618_t_to_slv(x : uint618_t) return std_logic_vector is
  variable rv : std_logic_vector(617 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint618_t(x : std_logic_vector) return uint618_t is
  variable rv : uint618_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int618_t_to_slv(x : int618_t) return std_logic_vector is
  variable rv : std_logic_vector(617 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int618_t(x : std_logic_vector) return int618_t is
  variable rv : int618_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint619_t_to_slv(x : uint619_t) return std_logic_vector is
  variable rv : std_logic_vector(618 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint619_t(x : std_logic_vector) return uint619_t is
  variable rv : uint619_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int619_t_to_slv(x : int619_t) return std_logic_vector is
  variable rv : std_logic_vector(618 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int619_t(x : std_logic_vector) return int619_t is
  variable rv : int619_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint620_t_to_slv(x : uint620_t) return std_logic_vector is
  variable rv : std_logic_vector(619 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint620_t(x : std_logic_vector) return uint620_t is
  variable rv : uint620_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int620_t_to_slv(x : int620_t) return std_logic_vector is
  variable rv : std_logic_vector(619 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int620_t(x : std_logic_vector) return int620_t is
  variable rv : int620_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint621_t_to_slv(x : uint621_t) return std_logic_vector is
  variable rv : std_logic_vector(620 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint621_t(x : std_logic_vector) return uint621_t is
  variable rv : uint621_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int621_t_to_slv(x : int621_t) return std_logic_vector is
  variable rv : std_logic_vector(620 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int621_t(x : std_logic_vector) return int621_t is
  variable rv : int621_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint622_t_to_slv(x : uint622_t) return std_logic_vector is
  variable rv : std_logic_vector(621 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint622_t(x : std_logic_vector) return uint622_t is
  variable rv : uint622_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int622_t_to_slv(x : int622_t) return std_logic_vector is
  variable rv : std_logic_vector(621 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int622_t(x : std_logic_vector) return int622_t is
  variable rv : int622_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint623_t_to_slv(x : uint623_t) return std_logic_vector is
  variable rv : std_logic_vector(622 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint623_t(x : std_logic_vector) return uint623_t is
  variable rv : uint623_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int623_t_to_slv(x : int623_t) return std_logic_vector is
  variable rv : std_logic_vector(622 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int623_t(x : std_logic_vector) return int623_t is
  variable rv : int623_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint624_t_to_slv(x : uint624_t) return std_logic_vector is
  variable rv : std_logic_vector(623 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint624_t(x : std_logic_vector) return uint624_t is
  variable rv : uint624_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int624_t_to_slv(x : int624_t) return std_logic_vector is
  variable rv : std_logic_vector(623 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int624_t(x : std_logic_vector) return int624_t is
  variable rv : int624_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint625_t_to_slv(x : uint625_t) return std_logic_vector is
  variable rv : std_logic_vector(624 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint625_t(x : std_logic_vector) return uint625_t is
  variable rv : uint625_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int625_t_to_slv(x : int625_t) return std_logic_vector is
  variable rv : std_logic_vector(624 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int625_t(x : std_logic_vector) return int625_t is
  variable rv : int625_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint626_t_to_slv(x : uint626_t) return std_logic_vector is
  variable rv : std_logic_vector(625 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint626_t(x : std_logic_vector) return uint626_t is
  variable rv : uint626_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int626_t_to_slv(x : int626_t) return std_logic_vector is
  variable rv : std_logic_vector(625 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int626_t(x : std_logic_vector) return int626_t is
  variable rv : int626_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint627_t_to_slv(x : uint627_t) return std_logic_vector is
  variable rv : std_logic_vector(626 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint627_t(x : std_logic_vector) return uint627_t is
  variable rv : uint627_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int627_t_to_slv(x : int627_t) return std_logic_vector is
  variable rv : std_logic_vector(626 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int627_t(x : std_logic_vector) return int627_t is
  variable rv : int627_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint628_t_to_slv(x : uint628_t) return std_logic_vector is
  variable rv : std_logic_vector(627 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint628_t(x : std_logic_vector) return uint628_t is
  variable rv : uint628_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int628_t_to_slv(x : int628_t) return std_logic_vector is
  variable rv : std_logic_vector(627 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int628_t(x : std_logic_vector) return int628_t is
  variable rv : int628_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint629_t_to_slv(x : uint629_t) return std_logic_vector is
  variable rv : std_logic_vector(628 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint629_t(x : std_logic_vector) return uint629_t is
  variable rv : uint629_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int629_t_to_slv(x : int629_t) return std_logic_vector is
  variable rv : std_logic_vector(628 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int629_t(x : std_logic_vector) return int629_t is
  variable rv : int629_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint630_t_to_slv(x : uint630_t) return std_logic_vector is
  variable rv : std_logic_vector(629 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint630_t(x : std_logic_vector) return uint630_t is
  variable rv : uint630_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int630_t_to_slv(x : int630_t) return std_logic_vector is
  variable rv : std_logic_vector(629 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int630_t(x : std_logic_vector) return int630_t is
  variable rv : int630_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint631_t_to_slv(x : uint631_t) return std_logic_vector is
  variable rv : std_logic_vector(630 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint631_t(x : std_logic_vector) return uint631_t is
  variable rv : uint631_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int631_t_to_slv(x : int631_t) return std_logic_vector is
  variable rv : std_logic_vector(630 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int631_t(x : std_logic_vector) return int631_t is
  variable rv : int631_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint632_t_to_slv(x : uint632_t) return std_logic_vector is
  variable rv : std_logic_vector(631 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint632_t(x : std_logic_vector) return uint632_t is
  variable rv : uint632_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int632_t_to_slv(x : int632_t) return std_logic_vector is
  variable rv : std_logic_vector(631 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int632_t(x : std_logic_vector) return int632_t is
  variable rv : int632_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint633_t_to_slv(x : uint633_t) return std_logic_vector is
  variable rv : std_logic_vector(632 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint633_t(x : std_logic_vector) return uint633_t is
  variable rv : uint633_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int633_t_to_slv(x : int633_t) return std_logic_vector is
  variable rv : std_logic_vector(632 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int633_t(x : std_logic_vector) return int633_t is
  variable rv : int633_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint634_t_to_slv(x : uint634_t) return std_logic_vector is
  variable rv : std_logic_vector(633 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint634_t(x : std_logic_vector) return uint634_t is
  variable rv : uint634_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int634_t_to_slv(x : int634_t) return std_logic_vector is
  variable rv : std_logic_vector(633 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int634_t(x : std_logic_vector) return int634_t is
  variable rv : int634_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint635_t_to_slv(x : uint635_t) return std_logic_vector is
  variable rv : std_logic_vector(634 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint635_t(x : std_logic_vector) return uint635_t is
  variable rv : uint635_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int635_t_to_slv(x : int635_t) return std_logic_vector is
  variable rv : std_logic_vector(634 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int635_t(x : std_logic_vector) return int635_t is
  variable rv : int635_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint636_t_to_slv(x : uint636_t) return std_logic_vector is
  variable rv : std_logic_vector(635 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint636_t(x : std_logic_vector) return uint636_t is
  variable rv : uint636_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int636_t_to_slv(x : int636_t) return std_logic_vector is
  variable rv : std_logic_vector(635 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int636_t(x : std_logic_vector) return int636_t is
  variable rv : int636_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint637_t_to_slv(x : uint637_t) return std_logic_vector is
  variable rv : std_logic_vector(636 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint637_t(x : std_logic_vector) return uint637_t is
  variable rv : uint637_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int637_t_to_slv(x : int637_t) return std_logic_vector is
  variable rv : std_logic_vector(636 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int637_t(x : std_logic_vector) return int637_t is
  variable rv : int637_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint638_t_to_slv(x : uint638_t) return std_logic_vector is
  variable rv : std_logic_vector(637 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint638_t(x : std_logic_vector) return uint638_t is
  variable rv : uint638_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int638_t_to_slv(x : int638_t) return std_logic_vector is
  variable rv : std_logic_vector(637 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int638_t(x : std_logic_vector) return int638_t is
  variable rv : int638_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint639_t_to_slv(x : uint639_t) return std_logic_vector is
  variable rv : std_logic_vector(638 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint639_t(x : std_logic_vector) return uint639_t is
  variable rv : uint639_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int639_t_to_slv(x : int639_t) return std_logic_vector is
  variable rv : std_logic_vector(638 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int639_t(x : std_logic_vector) return int639_t is
  variable rv : int639_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint640_t_to_slv(x : uint640_t) return std_logic_vector is
  variable rv : std_logic_vector(639 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint640_t(x : std_logic_vector) return uint640_t is
  variable rv : uint640_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int640_t_to_slv(x : int640_t) return std_logic_vector is
  variable rv : std_logic_vector(639 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int640_t(x : std_logic_vector) return int640_t is
  variable rv : int640_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint641_t_to_slv(x : uint641_t) return std_logic_vector is
  variable rv : std_logic_vector(640 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint641_t(x : std_logic_vector) return uint641_t is
  variable rv : uint641_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int641_t_to_slv(x : int641_t) return std_logic_vector is
  variable rv : std_logic_vector(640 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int641_t(x : std_logic_vector) return int641_t is
  variable rv : int641_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint642_t_to_slv(x : uint642_t) return std_logic_vector is
  variable rv : std_logic_vector(641 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint642_t(x : std_logic_vector) return uint642_t is
  variable rv : uint642_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int642_t_to_slv(x : int642_t) return std_logic_vector is
  variable rv : std_logic_vector(641 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int642_t(x : std_logic_vector) return int642_t is
  variable rv : int642_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint643_t_to_slv(x : uint643_t) return std_logic_vector is
  variable rv : std_logic_vector(642 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint643_t(x : std_logic_vector) return uint643_t is
  variable rv : uint643_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int643_t_to_slv(x : int643_t) return std_logic_vector is
  variable rv : std_logic_vector(642 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int643_t(x : std_logic_vector) return int643_t is
  variable rv : int643_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint644_t_to_slv(x : uint644_t) return std_logic_vector is
  variable rv : std_logic_vector(643 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint644_t(x : std_logic_vector) return uint644_t is
  variable rv : uint644_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int644_t_to_slv(x : int644_t) return std_logic_vector is
  variable rv : std_logic_vector(643 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int644_t(x : std_logic_vector) return int644_t is
  variable rv : int644_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint645_t_to_slv(x : uint645_t) return std_logic_vector is
  variable rv : std_logic_vector(644 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint645_t(x : std_logic_vector) return uint645_t is
  variable rv : uint645_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int645_t_to_slv(x : int645_t) return std_logic_vector is
  variable rv : std_logic_vector(644 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int645_t(x : std_logic_vector) return int645_t is
  variable rv : int645_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint646_t_to_slv(x : uint646_t) return std_logic_vector is
  variable rv : std_logic_vector(645 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint646_t(x : std_logic_vector) return uint646_t is
  variable rv : uint646_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int646_t_to_slv(x : int646_t) return std_logic_vector is
  variable rv : std_logic_vector(645 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int646_t(x : std_logic_vector) return int646_t is
  variable rv : int646_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint647_t_to_slv(x : uint647_t) return std_logic_vector is
  variable rv : std_logic_vector(646 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint647_t(x : std_logic_vector) return uint647_t is
  variable rv : uint647_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int647_t_to_slv(x : int647_t) return std_logic_vector is
  variable rv : std_logic_vector(646 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int647_t(x : std_logic_vector) return int647_t is
  variable rv : int647_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint648_t_to_slv(x : uint648_t) return std_logic_vector is
  variable rv : std_logic_vector(647 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint648_t(x : std_logic_vector) return uint648_t is
  variable rv : uint648_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int648_t_to_slv(x : int648_t) return std_logic_vector is
  variable rv : std_logic_vector(647 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int648_t(x : std_logic_vector) return int648_t is
  variable rv : int648_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint649_t_to_slv(x : uint649_t) return std_logic_vector is
  variable rv : std_logic_vector(648 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint649_t(x : std_logic_vector) return uint649_t is
  variable rv : uint649_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int649_t_to_slv(x : int649_t) return std_logic_vector is
  variable rv : std_logic_vector(648 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int649_t(x : std_logic_vector) return int649_t is
  variable rv : int649_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint650_t_to_slv(x : uint650_t) return std_logic_vector is
  variable rv : std_logic_vector(649 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint650_t(x : std_logic_vector) return uint650_t is
  variable rv : uint650_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int650_t_to_slv(x : int650_t) return std_logic_vector is
  variable rv : std_logic_vector(649 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int650_t(x : std_logic_vector) return int650_t is
  variable rv : int650_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint651_t_to_slv(x : uint651_t) return std_logic_vector is
  variable rv : std_logic_vector(650 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint651_t(x : std_logic_vector) return uint651_t is
  variable rv : uint651_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int651_t_to_slv(x : int651_t) return std_logic_vector is
  variable rv : std_logic_vector(650 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int651_t(x : std_logic_vector) return int651_t is
  variable rv : int651_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint652_t_to_slv(x : uint652_t) return std_logic_vector is
  variable rv : std_logic_vector(651 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint652_t(x : std_logic_vector) return uint652_t is
  variable rv : uint652_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int652_t_to_slv(x : int652_t) return std_logic_vector is
  variable rv : std_logic_vector(651 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int652_t(x : std_logic_vector) return int652_t is
  variable rv : int652_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint653_t_to_slv(x : uint653_t) return std_logic_vector is
  variable rv : std_logic_vector(652 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint653_t(x : std_logic_vector) return uint653_t is
  variable rv : uint653_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int653_t_to_slv(x : int653_t) return std_logic_vector is
  variable rv : std_logic_vector(652 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int653_t(x : std_logic_vector) return int653_t is
  variable rv : int653_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint654_t_to_slv(x : uint654_t) return std_logic_vector is
  variable rv : std_logic_vector(653 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint654_t(x : std_logic_vector) return uint654_t is
  variable rv : uint654_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int654_t_to_slv(x : int654_t) return std_logic_vector is
  variable rv : std_logic_vector(653 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int654_t(x : std_logic_vector) return int654_t is
  variable rv : int654_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint655_t_to_slv(x : uint655_t) return std_logic_vector is
  variable rv : std_logic_vector(654 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint655_t(x : std_logic_vector) return uint655_t is
  variable rv : uint655_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int655_t_to_slv(x : int655_t) return std_logic_vector is
  variable rv : std_logic_vector(654 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int655_t(x : std_logic_vector) return int655_t is
  variable rv : int655_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint656_t_to_slv(x : uint656_t) return std_logic_vector is
  variable rv : std_logic_vector(655 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint656_t(x : std_logic_vector) return uint656_t is
  variable rv : uint656_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int656_t_to_slv(x : int656_t) return std_logic_vector is
  variable rv : std_logic_vector(655 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int656_t(x : std_logic_vector) return int656_t is
  variable rv : int656_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint657_t_to_slv(x : uint657_t) return std_logic_vector is
  variable rv : std_logic_vector(656 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint657_t(x : std_logic_vector) return uint657_t is
  variable rv : uint657_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int657_t_to_slv(x : int657_t) return std_logic_vector is
  variable rv : std_logic_vector(656 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int657_t(x : std_logic_vector) return int657_t is
  variable rv : int657_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint658_t_to_slv(x : uint658_t) return std_logic_vector is
  variable rv : std_logic_vector(657 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint658_t(x : std_logic_vector) return uint658_t is
  variable rv : uint658_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int658_t_to_slv(x : int658_t) return std_logic_vector is
  variable rv : std_logic_vector(657 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int658_t(x : std_logic_vector) return int658_t is
  variable rv : int658_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint659_t_to_slv(x : uint659_t) return std_logic_vector is
  variable rv : std_logic_vector(658 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint659_t(x : std_logic_vector) return uint659_t is
  variable rv : uint659_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int659_t_to_slv(x : int659_t) return std_logic_vector is
  variable rv : std_logic_vector(658 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int659_t(x : std_logic_vector) return int659_t is
  variable rv : int659_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint660_t_to_slv(x : uint660_t) return std_logic_vector is
  variable rv : std_logic_vector(659 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint660_t(x : std_logic_vector) return uint660_t is
  variable rv : uint660_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int660_t_to_slv(x : int660_t) return std_logic_vector is
  variable rv : std_logic_vector(659 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int660_t(x : std_logic_vector) return int660_t is
  variable rv : int660_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint661_t_to_slv(x : uint661_t) return std_logic_vector is
  variable rv : std_logic_vector(660 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint661_t(x : std_logic_vector) return uint661_t is
  variable rv : uint661_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int661_t_to_slv(x : int661_t) return std_logic_vector is
  variable rv : std_logic_vector(660 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int661_t(x : std_logic_vector) return int661_t is
  variable rv : int661_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint662_t_to_slv(x : uint662_t) return std_logic_vector is
  variable rv : std_logic_vector(661 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint662_t(x : std_logic_vector) return uint662_t is
  variable rv : uint662_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int662_t_to_slv(x : int662_t) return std_logic_vector is
  variable rv : std_logic_vector(661 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int662_t(x : std_logic_vector) return int662_t is
  variable rv : int662_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint663_t_to_slv(x : uint663_t) return std_logic_vector is
  variable rv : std_logic_vector(662 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint663_t(x : std_logic_vector) return uint663_t is
  variable rv : uint663_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int663_t_to_slv(x : int663_t) return std_logic_vector is
  variable rv : std_logic_vector(662 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int663_t(x : std_logic_vector) return int663_t is
  variable rv : int663_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint664_t_to_slv(x : uint664_t) return std_logic_vector is
  variable rv : std_logic_vector(663 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint664_t(x : std_logic_vector) return uint664_t is
  variable rv : uint664_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int664_t_to_slv(x : int664_t) return std_logic_vector is
  variable rv : std_logic_vector(663 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int664_t(x : std_logic_vector) return int664_t is
  variable rv : int664_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint665_t_to_slv(x : uint665_t) return std_logic_vector is
  variable rv : std_logic_vector(664 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint665_t(x : std_logic_vector) return uint665_t is
  variable rv : uint665_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int665_t_to_slv(x : int665_t) return std_logic_vector is
  variable rv : std_logic_vector(664 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int665_t(x : std_logic_vector) return int665_t is
  variable rv : int665_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint666_t_to_slv(x : uint666_t) return std_logic_vector is
  variable rv : std_logic_vector(665 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint666_t(x : std_logic_vector) return uint666_t is
  variable rv : uint666_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int666_t_to_slv(x : int666_t) return std_logic_vector is
  variable rv : std_logic_vector(665 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int666_t(x : std_logic_vector) return int666_t is
  variable rv : int666_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint667_t_to_slv(x : uint667_t) return std_logic_vector is
  variable rv : std_logic_vector(666 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint667_t(x : std_logic_vector) return uint667_t is
  variable rv : uint667_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int667_t_to_slv(x : int667_t) return std_logic_vector is
  variable rv : std_logic_vector(666 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int667_t(x : std_logic_vector) return int667_t is
  variable rv : int667_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint668_t_to_slv(x : uint668_t) return std_logic_vector is
  variable rv : std_logic_vector(667 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint668_t(x : std_logic_vector) return uint668_t is
  variable rv : uint668_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int668_t_to_slv(x : int668_t) return std_logic_vector is
  variable rv : std_logic_vector(667 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int668_t(x : std_logic_vector) return int668_t is
  variable rv : int668_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint669_t_to_slv(x : uint669_t) return std_logic_vector is
  variable rv : std_logic_vector(668 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint669_t(x : std_logic_vector) return uint669_t is
  variable rv : uint669_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int669_t_to_slv(x : int669_t) return std_logic_vector is
  variable rv : std_logic_vector(668 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int669_t(x : std_logic_vector) return int669_t is
  variable rv : int669_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint670_t_to_slv(x : uint670_t) return std_logic_vector is
  variable rv : std_logic_vector(669 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint670_t(x : std_logic_vector) return uint670_t is
  variable rv : uint670_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int670_t_to_slv(x : int670_t) return std_logic_vector is
  variable rv : std_logic_vector(669 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int670_t(x : std_logic_vector) return int670_t is
  variable rv : int670_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint671_t_to_slv(x : uint671_t) return std_logic_vector is
  variable rv : std_logic_vector(670 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint671_t(x : std_logic_vector) return uint671_t is
  variable rv : uint671_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int671_t_to_slv(x : int671_t) return std_logic_vector is
  variable rv : std_logic_vector(670 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int671_t(x : std_logic_vector) return int671_t is
  variable rv : int671_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint672_t_to_slv(x : uint672_t) return std_logic_vector is
  variable rv : std_logic_vector(671 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint672_t(x : std_logic_vector) return uint672_t is
  variable rv : uint672_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int672_t_to_slv(x : int672_t) return std_logic_vector is
  variable rv : std_logic_vector(671 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int672_t(x : std_logic_vector) return int672_t is
  variable rv : int672_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint673_t_to_slv(x : uint673_t) return std_logic_vector is
  variable rv : std_logic_vector(672 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint673_t(x : std_logic_vector) return uint673_t is
  variable rv : uint673_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int673_t_to_slv(x : int673_t) return std_logic_vector is
  variable rv : std_logic_vector(672 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int673_t(x : std_logic_vector) return int673_t is
  variable rv : int673_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint674_t_to_slv(x : uint674_t) return std_logic_vector is
  variable rv : std_logic_vector(673 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint674_t(x : std_logic_vector) return uint674_t is
  variable rv : uint674_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int674_t_to_slv(x : int674_t) return std_logic_vector is
  variable rv : std_logic_vector(673 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int674_t(x : std_logic_vector) return int674_t is
  variable rv : int674_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint675_t_to_slv(x : uint675_t) return std_logic_vector is
  variable rv : std_logic_vector(674 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint675_t(x : std_logic_vector) return uint675_t is
  variable rv : uint675_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int675_t_to_slv(x : int675_t) return std_logic_vector is
  variable rv : std_logic_vector(674 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int675_t(x : std_logic_vector) return int675_t is
  variable rv : int675_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint676_t_to_slv(x : uint676_t) return std_logic_vector is
  variable rv : std_logic_vector(675 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint676_t(x : std_logic_vector) return uint676_t is
  variable rv : uint676_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int676_t_to_slv(x : int676_t) return std_logic_vector is
  variable rv : std_logic_vector(675 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int676_t(x : std_logic_vector) return int676_t is
  variable rv : int676_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint677_t_to_slv(x : uint677_t) return std_logic_vector is
  variable rv : std_logic_vector(676 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint677_t(x : std_logic_vector) return uint677_t is
  variable rv : uint677_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int677_t_to_slv(x : int677_t) return std_logic_vector is
  variable rv : std_logic_vector(676 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int677_t(x : std_logic_vector) return int677_t is
  variable rv : int677_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint678_t_to_slv(x : uint678_t) return std_logic_vector is
  variable rv : std_logic_vector(677 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint678_t(x : std_logic_vector) return uint678_t is
  variable rv : uint678_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int678_t_to_slv(x : int678_t) return std_logic_vector is
  variable rv : std_logic_vector(677 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int678_t(x : std_logic_vector) return int678_t is
  variable rv : int678_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint679_t_to_slv(x : uint679_t) return std_logic_vector is
  variable rv : std_logic_vector(678 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint679_t(x : std_logic_vector) return uint679_t is
  variable rv : uint679_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int679_t_to_slv(x : int679_t) return std_logic_vector is
  variable rv : std_logic_vector(678 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int679_t(x : std_logic_vector) return int679_t is
  variable rv : int679_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint680_t_to_slv(x : uint680_t) return std_logic_vector is
  variable rv : std_logic_vector(679 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint680_t(x : std_logic_vector) return uint680_t is
  variable rv : uint680_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int680_t_to_slv(x : int680_t) return std_logic_vector is
  variable rv : std_logic_vector(679 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int680_t(x : std_logic_vector) return int680_t is
  variable rv : int680_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint681_t_to_slv(x : uint681_t) return std_logic_vector is
  variable rv : std_logic_vector(680 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint681_t(x : std_logic_vector) return uint681_t is
  variable rv : uint681_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int681_t_to_slv(x : int681_t) return std_logic_vector is
  variable rv : std_logic_vector(680 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int681_t(x : std_logic_vector) return int681_t is
  variable rv : int681_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint682_t_to_slv(x : uint682_t) return std_logic_vector is
  variable rv : std_logic_vector(681 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint682_t(x : std_logic_vector) return uint682_t is
  variable rv : uint682_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int682_t_to_slv(x : int682_t) return std_logic_vector is
  variable rv : std_logic_vector(681 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int682_t(x : std_logic_vector) return int682_t is
  variable rv : int682_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint683_t_to_slv(x : uint683_t) return std_logic_vector is
  variable rv : std_logic_vector(682 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint683_t(x : std_logic_vector) return uint683_t is
  variable rv : uint683_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int683_t_to_slv(x : int683_t) return std_logic_vector is
  variable rv : std_logic_vector(682 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int683_t(x : std_logic_vector) return int683_t is
  variable rv : int683_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint684_t_to_slv(x : uint684_t) return std_logic_vector is
  variable rv : std_logic_vector(683 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint684_t(x : std_logic_vector) return uint684_t is
  variable rv : uint684_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int684_t_to_slv(x : int684_t) return std_logic_vector is
  variable rv : std_logic_vector(683 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int684_t(x : std_logic_vector) return int684_t is
  variable rv : int684_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint685_t_to_slv(x : uint685_t) return std_logic_vector is
  variable rv : std_logic_vector(684 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint685_t(x : std_logic_vector) return uint685_t is
  variable rv : uint685_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int685_t_to_slv(x : int685_t) return std_logic_vector is
  variable rv : std_logic_vector(684 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int685_t(x : std_logic_vector) return int685_t is
  variable rv : int685_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint686_t_to_slv(x : uint686_t) return std_logic_vector is
  variable rv : std_logic_vector(685 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint686_t(x : std_logic_vector) return uint686_t is
  variable rv : uint686_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int686_t_to_slv(x : int686_t) return std_logic_vector is
  variable rv : std_logic_vector(685 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int686_t(x : std_logic_vector) return int686_t is
  variable rv : int686_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint687_t_to_slv(x : uint687_t) return std_logic_vector is
  variable rv : std_logic_vector(686 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint687_t(x : std_logic_vector) return uint687_t is
  variable rv : uint687_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int687_t_to_slv(x : int687_t) return std_logic_vector is
  variable rv : std_logic_vector(686 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int687_t(x : std_logic_vector) return int687_t is
  variable rv : int687_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint688_t_to_slv(x : uint688_t) return std_logic_vector is
  variable rv : std_logic_vector(687 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint688_t(x : std_logic_vector) return uint688_t is
  variable rv : uint688_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int688_t_to_slv(x : int688_t) return std_logic_vector is
  variable rv : std_logic_vector(687 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int688_t(x : std_logic_vector) return int688_t is
  variable rv : int688_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint689_t_to_slv(x : uint689_t) return std_logic_vector is
  variable rv : std_logic_vector(688 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint689_t(x : std_logic_vector) return uint689_t is
  variable rv : uint689_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int689_t_to_slv(x : int689_t) return std_logic_vector is
  variable rv : std_logic_vector(688 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int689_t(x : std_logic_vector) return int689_t is
  variable rv : int689_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint690_t_to_slv(x : uint690_t) return std_logic_vector is
  variable rv : std_logic_vector(689 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint690_t(x : std_logic_vector) return uint690_t is
  variable rv : uint690_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int690_t_to_slv(x : int690_t) return std_logic_vector is
  variable rv : std_logic_vector(689 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int690_t(x : std_logic_vector) return int690_t is
  variable rv : int690_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint691_t_to_slv(x : uint691_t) return std_logic_vector is
  variable rv : std_logic_vector(690 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint691_t(x : std_logic_vector) return uint691_t is
  variable rv : uint691_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int691_t_to_slv(x : int691_t) return std_logic_vector is
  variable rv : std_logic_vector(690 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int691_t(x : std_logic_vector) return int691_t is
  variable rv : int691_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint692_t_to_slv(x : uint692_t) return std_logic_vector is
  variable rv : std_logic_vector(691 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint692_t(x : std_logic_vector) return uint692_t is
  variable rv : uint692_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int692_t_to_slv(x : int692_t) return std_logic_vector is
  variable rv : std_logic_vector(691 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int692_t(x : std_logic_vector) return int692_t is
  variable rv : int692_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint693_t_to_slv(x : uint693_t) return std_logic_vector is
  variable rv : std_logic_vector(692 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint693_t(x : std_logic_vector) return uint693_t is
  variable rv : uint693_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int693_t_to_slv(x : int693_t) return std_logic_vector is
  variable rv : std_logic_vector(692 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int693_t(x : std_logic_vector) return int693_t is
  variable rv : int693_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint694_t_to_slv(x : uint694_t) return std_logic_vector is
  variable rv : std_logic_vector(693 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint694_t(x : std_logic_vector) return uint694_t is
  variable rv : uint694_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int694_t_to_slv(x : int694_t) return std_logic_vector is
  variable rv : std_logic_vector(693 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int694_t(x : std_logic_vector) return int694_t is
  variable rv : int694_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint695_t_to_slv(x : uint695_t) return std_logic_vector is
  variable rv : std_logic_vector(694 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint695_t(x : std_logic_vector) return uint695_t is
  variable rv : uint695_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int695_t_to_slv(x : int695_t) return std_logic_vector is
  variable rv : std_logic_vector(694 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int695_t(x : std_logic_vector) return int695_t is
  variable rv : int695_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint696_t_to_slv(x : uint696_t) return std_logic_vector is
  variable rv : std_logic_vector(695 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint696_t(x : std_logic_vector) return uint696_t is
  variable rv : uint696_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int696_t_to_slv(x : int696_t) return std_logic_vector is
  variable rv : std_logic_vector(695 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int696_t(x : std_logic_vector) return int696_t is
  variable rv : int696_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint697_t_to_slv(x : uint697_t) return std_logic_vector is
  variable rv : std_logic_vector(696 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint697_t(x : std_logic_vector) return uint697_t is
  variable rv : uint697_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int697_t_to_slv(x : int697_t) return std_logic_vector is
  variable rv : std_logic_vector(696 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int697_t(x : std_logic_vector) return int697_t is
  variable rv : int697_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint698_t_to_slv(x : uint698_t) return std_logic_vector is
  variable rv : std_logic_vector(697 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint698_t(x : std_logic_vector) return uint698_t is
  variable rv : uint698_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int698_t_to_slv(x : int698_t) return std_logic_vector is
  variable rv : std_logic_vector(697 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int698_t(x : std_logic_vector) return int698_t is
  variable rv : int698_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint699_t_to_slv(x : uint699_t) return std_logic_vector is
  variable rv : std_logic_vector(698 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint699_t(x : std_logic_vector) return uint699_t is
  variable rv : uint699_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int699_t_to_slv(x : int699_t) return std_logic_vector is
  variable rv : std_logic_vector(698 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int699_t(x : std_logic_vector) return int699_t is
  variable rv : int699_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint700_t_to_slv(x : uint700_t) return std_logic_vector is
  variable rv : std_logic_vector(699 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint700_t(x : std_logic_vector) return uint700_t is
  variable rv : uint700_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int700_t_to_slv(x : int700_t) return std_logic_vector is
  variable rv : std_logic_vector(699 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int700_t(x : std_logic_vector) return int700_t is
  variable rv : int700_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint701_t_to_slv(x : uint701_t) return std_logic_vector is
  variable rv : std_logic_vector(700 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint701_t(x : std_logic_vector) return uint701_t is
  variable rv : uint701_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int701_t_to_slv(x : int701_t) return std_logic_vector is
  variable rv : std_logic_vector(700 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int701_t(x : std_logic_vector) return int701_t is
  variable rv : int701_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint702_t_to_slv(x : uint702_t) return std_logic_vector is
  variable rv : std_logic_vector(701 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint702_t(x : std_logic_vector) return uint702_t is
  variable rv : uint702_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int702_t_to_slv(x : int702_t) return std_logic_vector is
  variable rv : std_logic_vector(701 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int702_t(x : std_logic_vector) return int702_t is
  variable rv : int702_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint703_t_to_slv(x : uint703_t) return std_logic_vector is
  variable rv : std_logic_vector(702 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint703_t(x : std_logic_vector) return uint703_t is
  variable rv : uint703_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int703_t_to_slv(x : int703_t) return std_logic_vector is
  variable rv : std_logic_vector(702 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int703_t(x : std_logic_vector) return int703_t is
  variable rv : int703_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint704_t_to_slv(x : uint704_t) return std_logic_vector is
  variable rv : std_logic_vector(703 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint704_t(x : std_logic_vector) return uint704_t is
  variable rv : uint704_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int704_t_to_slv(x : int704_t) return std_logic_vector is
  variable rv : std_logic_vector(703 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int704_t(x : std_logic_vector) return int704_t is
  variable rv : int704_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint705_t_to_slv(x : uint705_t) return std_logic_vector is
  variable rv : std_logic_vector(704 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint705_t(x : std_logic_vector) return uint705_t is
  variable rv : uint705_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int705_t_to_slv(x : int705_t) return std_logic_vector is
  variable rv : std_logic_vector(704 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int705_t(x : std_logic_vector) return int705_t is
  variable rv : int705_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint706_t_to_slv(x : uint706_t) return std_logic_vector is
  variable rv : std_logic_vector(705 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint706_t(x : std_logic_vector) return uint706_t is
  variable rv : uint706_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int706_t_to_slv(x : int706_t) return std_logic_vector is
  variable rv : std_logic_vector(705 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int706_t(x : std_logic_vector) return int706_t is
  variable rv : int706_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint707_t_to_slv(x : uint707_t) return std_logic_vector is
  variable rv : std_logic_vector(706 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint707_t(x : std_logic_vector) return uint707_t is
  variable rv : uint707_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int707_t_to_slv(x : int707_t) return std_logic_vector is
  variable rv : std_logic_vector(706 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int707_t(x : std_logic_vector) return int707_t is
  variable rv : int707_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint708_t_to_slv(x : uint708_t) return std_logic_vector is
  variable rv : std_logic_vector(707 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint708_t(x : std_logic_vector) return uint708_t is
  variable rv : uint708_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int708_t_to_slv(x : int708_t) return std_logic_vector is
  variable rv : std_logic_vector(707 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int708_t(x : std_logic_vector) return int708_t is
  variable rv : int708_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint709_t_to_slv(x : uint709_t) return std_logic_vector is
  variable rv : std_logic_vector(708 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint709_t(x : std_logic_vector) return uint709_t is
  variable rv : uint709_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int709_t_to_slv(x : int709_t) return std_logic_vector is
  variable rv : std_logic_vector(708 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int709_t(x : std_logic_vector) return int709_t is
  variable rv : int709_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint710_t_to_slv(x : uint710_t) return std_logic_vector is
  variable rv : std_logic_vector(709 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint710_t(x : std_logic_vector) return uint710_t is
  variable rv : uint710_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int710_t_to_slv(x : int710_t) return std_logic_vector is
  variable rv : std_logic_vector(709 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int710_t(x : std_logic_vector) return int710_t is
  variable rv : int710_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint711_t_to_slv(x : uint711_t) return std_logic_vector is
  variable rv : std_logic_vector(710 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint711_t(x : std_logic_vector) return uint711_t is
  variable rv : uint711_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int711_t_to_slv(x : int711_t) return std_logic_vector is
  variable rv : std_logic_vector(710 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int711_t(x : std_logic_vector) return int711_t is
  variable rv : int711_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint712_t_to_slv(x : uint712_t) return std_logic_vector is
  variable rv : std_logic_vector(711 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint712_t(x : std_logic_vector) return uint712_t is
  variable rv : uint712_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int712_t_to_slv(x : int712_t) return std_logic_vector is
  variable rv : std_logic_vector(711 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int712_t(x : std_logic_vector) return int712_t is
  variable rv : int712_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint713_t_to_slv(x : uint713_t) return std_logic_vector is
  variable rv : std_logic_vector(712 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint713_t(x : std_logic_vector) return uint713_t is
  variable rv : uint713_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int713_t_to_slv(x : int713_t) return std_logic_vector is
  variable rv : std_logic_vector(712 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int713_t(x : std_logic_vector) return int713_t is
  variable rv : int713_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint714_t_to_slv(x : uint714_t) return std_logic_vector is
  variable rv : std_logic_vector(713 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint714_t(x : std_logic_vector) return uint714_t is
  variable rv : uint714_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int714_t_to_slv(x : int714_t) return std_logic_vector is
  variable rv : std_logic_vector(713 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int714_t(x : std_logic_vector) return int714_t is
  variable rv : int714_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint715_t_to_slv(x : uint715_t) return std_logic_vector is
  variable rv : std_logic_vector(714 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint715_t(x : std_logic_vector) return uint715_t is
  variable rv : uint715_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int715_t_to_slv(x : int715_t) return std_logic_vector is
  variable rv : std_logic_vector(714 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int715_t(x : std_logic_vector) return int715_t is
  variable rv : int715_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint716_t_to_slv(x : uint716_t) return std_logic_vector is
  variable rv : std_logic_vector(715 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint716_t(x : std_logic_vector) return uint716_t is
  variable rv : uint716_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int716_t_to_slv(x : int716_t) return std_logic_vector is
  variable rv : std_logic_vector(715 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int716_t(x : std_logic_vector) return int716_t is
  variable rv : int716_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint717_t_to_slv(x : uint717_t) return std_logic_vector is
  variable rv : std_logic_vector(716 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint717_t(x : std_logic_vector) return uint717_t is
  variable rv : uint717_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int717_t_to_slv(x : int717_t) return std_logic_vector is
  variable rv : std_logic_vector(716 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int717_t(x : std_logic_vector) return int717_t is
  variable rv : int717_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint718_t_to_slv(x : uint718_t) return std_logic_vector is
  variable rv : std_logic_vector(717 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint718_t(x : std_logic_vector) return uint718_t is
  variable rv : uint718_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int718_t_to_slv(x : int718_t) return std_logic_vector is
  variable rv : std_logic_vector(717 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int718_t(x : std_logic_vector) return int718_t is
  variable rv : int718_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint719_t_to_slv(x : uint719_t) return std_logic_vector is
  variable rv : std_logic_vector(718 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint719_t(x : std_logic_vector) return uint719_t is
  variable rv : uint719_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int719_t_to_slv(x : int719_t) return std_logic_vector is
  variable rv : std_logic_vector(718 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int719_t(x : std_logic_vector) return int719_t is
  variable rv : int719_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint720_t_to_slv(x : uint720_t) return std_logic_vector is
  variable rv : std_logic_vector(719 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint720_t(x : std_logic_vector) return uint720_t is
  variable rv : uint720_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int720_t_to_slv(x : int720_t) return std_logic_vector is
  variable rv : std_logic_vector(719 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int720_t(x : std_logic_vector) return int720_t is
  variable rv : int720_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint721_t_to_slv(x : uint721_t) return std_logic_vector is
  variable rv : std_logic_vector(720 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint721_t(x : std_logic_vector) return uint721_t is
  variable rv : uint721_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int721_t_to_slv(x : int721_t) return std_logic_vector is
  variable rv : std_logic_vector(720 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int721_t(x : std_logic_vector) return int721_t is
  variable rv : int721_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint722_t_to_slv(x : uint722_t) return std_logic_vector is
  variable rv : std_logic_vector(721 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint722_t(x : std_logic_vector) return uint722_t is
  variable rv : uint722_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int722_t_to_slv(x : int722_t) return std_logic_vector is
  variable rv : std_logic_vector(721 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int722_t(x : std_logic_vector) return int722_t is
  variable rv : int722_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint723_t_to_slv(x : uint723_t) return std_logic_vector is
  variable rv : std_logic_vector(722 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint723_t(x : std_logic_vector) return uint723_t is
  variable rv : uint723_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int723_t_to_slv(x : int723_t) return std_logic_vector is
  variable rv : std_logic_vector(722 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int723_t(x : std_logic_vector) return int723_t is
  variable rv : int723_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint724_t_to_slv(x : uint724_t) return std_logic_vector is
  variable rv : std_logic_vector(723 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint724_t(x : std_logic_vector) return uint724_t is
  variable rv : uint724_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int724_t_to_slv(x : int724_t) return std_logic_vector is
  variable rv : std_logic_vector(723 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int724_t(x : std_logic_vector) return int724_t is
  variable rv : int724_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint725_t_to_slv(x : uint725_t) return std_logic_vector is
  variable rv : std_logic_vector(724 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint725_t(x : std_logic_vector) return uint725_t is
  variable rv : uint725_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int725_t_to_slv(x : int725_t) return std_logic_vector is
  variable rv : std_logic_vector(724 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int725_t(x : std_logic_vector) return int725_t is
  variable rv : int725_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint726_t_to_slv(x : uint726_t) return std_logic_vector is
  variable rv : std_logic_vector(725 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint726_t(x : std_logic_vector) return uint726_t is
  variable rv : uint726_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int726_t_to_slv(x : int726_t) return std_logic_vector is
  variable rv : std_logic_vector(725 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int726_t(x : std_logic_vector) return int726_t is
  variable rv : int726_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint727_t_to_slv(x : uint727_t) return std_logic_vector is
  variable rv : std_logic_vector(726 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint727_t(x : std_logic_vector) return uint727_t is
  variable rv : uint727_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int727_t_to_slv(x : int727_t) return std_logic_vector is
  variable rv : std_logic_vector(726 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int727_t(x : std_logic_vector) return int727_t is
  variable rv : int727_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint728_t_to_slv(x : uint728_t) return std_logic_vector is
  variable rv : std_logic_vector(727 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint728_t(x : std_logic_vector) return uint728_t is
  variable rv : uint728_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int728_t_to_slv(x : int728_t) return std_logic_vector is
  variable rv : std_logic_vector(727 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int728_t(x : std_logic_vector) return int728_t is
  variable rv : int728_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint729_t_to_slv(x : uint729_t) return std_logic_vector is
  variable rv : std_logic_vector(728 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint729_t(x : std_logic_vector) return uint729_t is
  variable rv : uint729_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int729_t_to_slv(x : int729_t) return std_logic_vector is
  variable rv : std_logic_vector(728 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int729_t(x : std_logic_vector) return int729_t is
  variable rv : int729_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint730_t_to_slv(x : uint730_t) return std_logic_vector is
  variable rv : std_logic_vector(729 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint730_t(x : std_logic_vector) return uint730_t is
  variable rv : uint730_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int730_t_to_slv(x : int730_t) return std_logic_vector is
  variable rv : std_logic_vector(729 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int730_t(x : std_logic_vector) return int730_t is
  variable rv : int730_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint731_t_to_slv(x : uint731_t) return std_logic_vector is
  variable rv : std_logic_vector(730 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint731_t(x : std_logic_vector) return uint731_t is
  variable rv : uint731_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int731_t_to_slv(x : int731_t) return std_logic_vector is
  variable rv : std_logic_vector(730 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int731_t(x : std_logic_vector) return int731_t is
  variable rv : int731_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint732_t_to_slv(x : uint732_t) return std_logic_vector is
  variable rv : std_logic_vector(731 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint732_t(x : std_logic_vector) return uint732_t is
  variable rv : uint732_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int732_t_to_slv(x : int732_t) return std_logic_vector is
  variable rv : std_logic_vector(731 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int732_t(x : std_logic_vector) return int732_t is
  variable rv : int732_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint733_t_to_slv(x : uint733_t) return std_logic_vector is
  variable rv : std_logic_vector(732 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint733_t(x : std_logic_vector) return uint733_t is
  variable rv : uint733_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int733_t_to_slv(x : int733_t) return std_logic_vector is
  variable rv : std_logic_vector(732 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int733_t(x : std_logic_vector) return int733_t is
  variable rv : int733_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint734_t_to_slv(x : uint734_t) return std_logic_vector is
  variable rv : std_logic_vector(733 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint734_t(x : std_logic_vector) return uint734_t is
  variable rv : uint734_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int734_t_to_slv(x : int734_t) return std_logic_vector is
  variable rv : std_logic_vector(733 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int734_t(x : std_logic_vector) return int734_t is
  variable rv : int734_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint735_t_to_slv(x : uint735_t) return std_logic_vector is
  variable rv : std_logic_vector(734 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint735_t(x : std_logic_vector) return uint735_t is
  variable rv : uint735_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int735_t_to_slv(x : int735_t) return std_logic_vector is
  variable rv : std_logic_vector(734 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int735_t(x : std_logic_vector) return int735_t is
  variable rv : int735_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint736_t_to_slv(x : uint736_t) return std_logic_vector is
  variable rv : std_logic_vector(735 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint736_t(x : std_logic_vector) return uint736_t is
  variable rv : uint736_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int736_t_to_slv(x : int736_t) return std_logic_vector is
  variable rv : std_logic_vector(735 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int736_t(x : std_logic_vector) return int736_t is
  variable rv : int736_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint737_t_to_slv(x : uint737_t) return std_logic_vector is
  variable rv : std_logic_vector(736 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint737_t(x : std_logic_vector) return uint737_t is
  variable rv : uint737_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int737_t_to_slv(x : int737_t) return std_logic_vector is
  variable rv : std_logic_vector(736 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int737_t(x : std_logic_vector) return int737_t is
  variable rv : int737_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint738_t_to_slv(x : uint738_t) return std_logic_vector is
  variable rv : std_logic_vector(737 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint738_t(x : std_logic_vector) return uint738_t is
  variable rv : uint738_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int738_t_to_slv(x : int738_t) return std_logic_vector is
  variable rv : std_logic_vector(737 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int738_t(x : std_logic_vector) return int738_t is
  variable rv : int738_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint739_t_to_slv(x : uint739_t) return std_logic_vector is
  variable rv : std_logic_vector(738 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint739_t(x : std_logic_vector) return uint739_t is
  variable rv : uint739_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int739_t_to_slv(x : int739_t) return std_logic_vector is
  variable rv : std_logic_vector(738 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int739_t(x : std_logic_vector) return int739_t is
  variable rv : int739_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint740_t_to_slv(x : uint740_t) return std_logic_vector is
  variable rv : std_logic_vector(739 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint740_t(x : std_logic_vector) return uint740_t is
  variable rv : uint740_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int740_t_to_slv(x : int740_t) return std_logic_vector is
  variable rv : std_logic_vector(739 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int740_t(x : std_logic_vector) return int740_t is
  variable rv : int740_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint741_t_to_slv(x : uint741_t) return std_logic_vector is
  variable rv : std_logic_vector(740 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint741_t(x : std_logic_vector) return uint741_t is
  variable rv : uint741_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int741_t_to_slv(x : int741_t) return std_logic_vector is
  variable rv : std_logic_vector(740 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int741_t(x : std_logic_vector) return int741_t is
  variable rv : int741_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint742_t_to_slv(x : uint742_t) return std_logic_vector is
  variable rv : std_logic_vector(741 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint742_t(x : std_logic_vector) return uint742_t is
  variable rv : uint742_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int742_t_to_slv(x : int742_t) return std_logic_vector is
  variable rv : std_logic_vector(741 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int742_t(x : std_logic_vector) return int742_t is
  variable rv : int742_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint743_t_to_slv(x : uint743_t) return std_logic_vector is
  variable rv : std_logic_vector(742 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint743_t(x : std_logic_vector) return uint743_t is
  variable rv : uint743_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int743_t_to_slv(x : int743_t) return std_logic_vector is
  variable rv : std_logic_vector(742 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int743_t(x : std_logic_vector) return int743_t is
  variable rv : int743_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint744_t_to_slv(x : uint744_t) return std_logic_vector is
  variable rv : std_logic_vector(743 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint744_t(x : std_logic_vector) return uint744_t is
  variable rv : uint744_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int744_t_to_slv(x : int744_t) return std_logic_vector is
  variable rv : std_logic_vector(743 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int744_t(x : std_logic_vector) return int744_t is
  variable rv : int744_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint745_t_to_slv(x : uint745_t) return std_logic_vector is
  variable rv : std_logic_vector(744 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint745_t(x : std_logic_vector) return uint745_t is
  variable rv : uint745_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int745_t_to_slv(x : int745_t) return std_logic_vector is
  variable rv : std_logic_vector(744 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int745_t(x : std_logic_vector) return int745_t is
  variable rv : int745_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint746_t_to_slv(x : uint746_t) return std_logic_vector is
  variable rv : std_logic_vector(745 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint746_t(x : std_logic_vector) return uint746_t is
  variable rv : uint746_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int746_t_to_slv(x : int746_t) return std_logic_vector is
  variable rv : std_logic_vector(745 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int746_t(x : std_logic_vector) return int746_t is
  variable rv : int746_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint747_t_to_slv(x : uint747_t) return std_logic_vector is
  variable rv : std_logic_vector(746 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint747_t(x : std_logic_vector) return uint747_t is
  variable rv : uint747_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int747_t_to_slv(x : int747_t) return std_logic_vector is
  variable rv : std_logic_vector(746 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int747_t(x : std_logic_vector) return int747_t is
  variable rv : int747_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint748_t_to_slv(x : uint748_t) return std_logic_vector is
  variable rv : std_logic_vector(747 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint748_t(x : std_logic_vector) return uint748_t is
  variable rv : uint748_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int748_t_to_slv(x : int748_t) return std_logic_vector is
  variable rv : std_logic_vector(747 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int748_t(x : std_logic_vector) return int748_t is
  variable rv : int748_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint749_t_to_slv(x : uint749_t) return std_logic_vector is
  variable rv : std_logic_vector(748 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint749_t(x : std_logic_vector) return uint749_t is
  variable rv : uint749_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int749_t_to_slv(x : int749_t) return std_logic_vector is
  variable rv : std_logic_vector(748 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int749_t(x : std_logic_vector) return int749_t is
  variable rv : int749_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint750_t_to_slv(x : uint750_t) return std_logic_vector is
  variable rv : std_logic_vector(749 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint750_t(x : std_logic_vector) return uint750_t is
  variable rv : uint750_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int750_t_to_slv(x : int750_t) return std_logic_vector is
  variable rv : std_logic_vector(749 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int750_t(x : std_logic_vector) return int750_t is
  variable rv : int750_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint751_t_to_slv(x : uint751_t) return std_logic_vector is
  variable rv : std_logic_vector(750 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint751_t(x : std_logic_vector) return uint751_t is
  variable rv : uint751_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int751_t_to_slv(x : int751_t) return std_logic_vector is
  variable rv : std_logic_vector(750 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int751_t(x : std_logic_vector) return int751_t is
  variable rv : int751_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint752_t_to_slv(x : uint752_t) return std_logic_vector is
  variable rv : std_logic_vector(751 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint752_t(x : std_logic_vector) return uint752_t is
  variable rv : uint752_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int752_t_to_slv(x : int752_t) return std_logic_vector is
  variable rv : std_logic_vector(751 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int752_t(x : std_logic_vector) return int752_t is
  variable rv : int752_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint753_t_to_slv(x : uint753_t) return std_logic_vector is
  variable rv : std_logic_vector(752 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint753_t(x : std_logic_vector) return uint753_t is
  variable rv : uint753_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int753_t_to_slv(x : int753_t) return std_logic_vector is
  variable rv : std_logic_vector(752 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int753_t(x : std_logic_vector) return int753_t is
  variable rv : int753_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint754_t_to_slv(x : uint754_t) return std_logic_vector is
  variable rv : std_logic_vector(753 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint754_t(x : std_logic_vector) return uint754_t is
  variable rv : uint754_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int754_t_to_slv(x : int754_t) return std_logic_vector is
  variable rv : std_logic_vector(753 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int754_t(x : std_logic_vector) return int754_t is
  variable rv : int754_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint755_t_to_slv(x : uint755_t) return std_logic_vector is
  variable rv : std_logic_vector(754 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint755_t(x : std_logic_vector) return uint755_t is
  variable rv : uint755_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int755_t_to_slv(x : int755_t) return std_logic_vector is
  variable rv : std_logic_vector(754 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int755_t(x : std_logic_vector) return int755_t is
  variable rv : int755_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint756_t_to_slv(x : uint756_t) return std_logic_vector is
  variable rv : std_logic_vector(755 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint756_t(x : std_logic_vector) return uint756_t is
  variable rv : uint756_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int756_t_to_slv(x : int756_t) return std_logic_vector is
  variable rv : std_logic_vector(755 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int756_t(x : std_logic_vector) return int756_t is
  variable rv : int756_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint757_t_to_slv(x : uint757_t) return std_logic_vector is
  variable rv : std_logic_vector(756 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint757_t(x : std_logic_vector) return uint757_t is
  variable rv : uint757_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int757_t_to_slv(x : int757_t) return std_logic_vector is
  variable rv : std_logic_vector(756 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int757_t(x : std_logic_vector) return int757_t is
  variable rv : int757_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint758_t_to_slv(x : uint758_t) return std_logic_vector is
  variable rv : std_logic_vector(757 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint758_t(x : std_logic_vector) return uint758_t is
  variable rv : uint758_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int758_t_to_slv(x : int758_t) return std_logic_vector is
  variable rv : std_logic_vector(757 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int758_t(x : std_logic_vector) return int758_t is
  variable rv : int758_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint759_t_to_slv(x : uint759_t) return std_logic_vector is
  variable rv : std_logic_vector(758 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint759_t(x : std_logic_vector) return uint759_t is
  variable rv : uint759_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int759_t_to_slv(x : int759_t) return std_logic_vector is
  variable rv : std_logic_vector(758 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int759_t(x : std_logic_vector) return int759_t is
  variable rv : int759_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint760_t_to_slv(x : uint760_t) return std_logic_vector is
  variable rv : std_logic_vector(759 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint760_t(x : std_logic_vector) return uint760_t is
  variable rv : uint760_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int760_t_to_slv(x : int760_t) return std_logic_vector is
  variable rv : std_logic_vector(759 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int760_t(x : std_logic_vector) return int760_t is
  variable rv : int760_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint761_t_to_slv(x : uint761_t) return std_logic_vector is
  variable rv : std_logic_vector(760 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint761_t(x : std_logic_vector) return uint761_t is
  variable rv : uint761_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int761_t_to_slv(x : int761_t) return std_logic_vector is
  variable rv : std_logic_vector(760 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int761_t(x : std_logic_vector) return int761_t is
  variable rv : int761_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint762_t_to_slv(x : uint762_t) return std_logic_vector is
  variable rv : std_logic_vector(761 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint762_t(x : std_logic_vector) return uint762_t is
  variable rv : uint762_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int762_t_to_slv(x : int762_t) return std_logic_vector is
  variable rv : std_logic_vector(761 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int762_t(x : std_logic_vector) return int762_t is
  variable rv : int762_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint763_t_to_slv(x : uint763_t) return std_logic_vector is
  variable rv : std_logic_vector(762 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint763_t(x : std_logic_vector) return uint763_t is
  variable rv : uint763_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int763_t_to_slv(x : int763_t) return std_logic_vector is
  variable rv : std_logic_vector(762 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int763_t(x : std_logic_vector) return int763_t is
  variable rv : int763_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint764_t_to_slv(x : uint764_t) return std_logic_vector is
  variable rv : std_logic_vector(763 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint764_t(x : std_logic_vector) return uint764_t is
  variable rv : uint764_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int764_t_to_slv(x : int764_t) return std_logic_vector is
  variable rv : std_logic_vector(763 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int764_t(x : std_logic_vector) return int764_t is
  variable rv : int764_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint765_t_to_slv(x : uint765_t) return std_logic_vector is
  variable rv : std_logic_vector(764 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint765_t(x : std_logic_vector) return uint765_t is
  variable rv : uint765_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int765_t_to_slv(x : int765_t) return std_logic_vector is
  variable rv : std_logic_vector(764 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int765_t(x : std_logic_vector) return int765_t is
  variable rv : int765_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint766_t_to_slv(x : uint766_t) return std_logic_vector is
  variable rv : std_logic_vector(765 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint766_t(x : std_logic_vector) return uint766_t is
  variable rv : uint766_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int766_t_to_slv(x : int766_t) return std_logic_vector is
  variable rv : std_logic_vector(765 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int766_t(x : std_logic_vector) return int766_t is
  variable rv : int766_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint767_t_to_slv(x : uint767_t) return std_logic_vector is
  variable rv : std_logic_vector(766 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint767_t(x : std_logic_vector) return uint767_t is
  variable rv : uint767_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int767_t_to_slv(x : int767_t) return std_logic_vector is
  variable rv : std_logic_vector(766 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int767_t(x : std_logic_vector) return int767_t is
  variable rv : int767_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint768_t_to_slv(x : uint768_t) return std_logic_vector is
  variable rv : std_logic_vector(767 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint768_t(x : std_logic_vector) return uint768_t is
  variable rv : uint768_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int768_t_to_slv(x : int768_t) return std_logic_vector is
  variable rv : std_logic_vector(767 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int768_t(x : std_logic_vector) return int768_t is
  variable rv : int768_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint769_t_to_slv(x : uint769_t) return std_logic_vector is
  variable rv : std_logic_vector(768 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint769_t(x : std_logic_vector) return uint769_t is
  variable rv : uint769_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int769_t_to_slv(x : int769_t) return std_logic_vector is
  variable rv : std_logic_vector(768 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int769_t(x : std_logic_vector) return int769_t is
  variable rv : int769_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint770_t_to_slv(x : uint770_t) return std_logic_vector is
  variable rv : std_logic_vector(769 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint770_t(x : std_logic_vector) return uint770_t is
  variable rv : uint770_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int770_t_to_slv(x : int770_t) return std_logic_vector is
  variable rv : std_logic_vector(769 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int770_t(x : std_logic_vector) return int770_t is
  variable rv : int770_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint771_t_to_slv(x : uint771_t) return std_logic_vector is
  variable rv : std_logic_vector(770 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint771_t(x : std_logic_vector) return uint771_t is
  variable rv : uint771_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int771_t_to_slv(x : int771_t) return std_logic_vector is
  variable rv : std_logic_vector(770 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int771_t(x : std_logic_vector) return int771_t is
  variable rv : int771_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint772_t_to_slv(x : uint772_t) return std_logic_vector is
  variable rv : std_logic_vector(771 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint772_t(x : std_logic_vector) return uint772_t is
  variable rv : uint772_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int772_t_to_slv(x : int772_t) return std_logic_vector is
  variable rv : std_logic_vector(771 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int772_t(x : std_logic_vector) return int772_t is
  variable rv : int772_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint773_t_to_slv(x : uint773_t) return std_logic_vector is
  variable rv : std_logic_vector(772 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint773_t(x : std_logic_vector) return uint773_t is
  variable rv : uint773_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int773_t_to_slv(x : int773_t) return std_logic_vector is
  variable rv : std_logic_vector(772 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int773_t(x : std_logic_vector) return int773_t is
  variable rv : int773_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint774_t_to_slv(x : uint774_t) return std_logic_vector is
  variable rv : std_logic_vector(773 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint774_t(x : std_logic_vector) return uint774_t is
  variable rv : uint774_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int774_t_to_slv(x : int774_t) return std_logic_vector is
  variable rv : std_logic_vector(773 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int774_t(x : std_logic_vector) return int774_t is
  variable rv : int774_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint775_t_to_slv(x : uint775_t) return std_logic_vector is
  variable rv : std_logic_vector(774 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint775_t(x : std_logic_vector) return uint775_t is
  variable rv : uint775_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int775_t_to_slv(x : int775_t) return std_logic_vector is
  variable rv : std_logic_vector(774 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int775_t(x : std_logic_vector) return int775_t is
  variable rv : int775_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint776_t_to_slv(x : uint776_t) return std_logic_vector is
  variable rv : std_logic_vector(775 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint776_t(x : std_logic_vector) return uint776_t is
  variable rv : uint776_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int776_t_to_slv(x : int776_t) return std_logic_vector is
  variable rv : std_logic_vector(775 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int776_t(x : std_logic_vector) return int776_t is
  variable rv : int776_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint777_t_to_slv(x : uint777_t) return std_logic_vector is
  variable rv : std_logic_vector(776 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint777_t(x : std_logic_vector) return uint777_t is
  variable rv : uint777_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int777_t_to_slv(x : int777_t) return std_logic_vector is
  variable rv : std_logic_vector(776 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int777_t(x : std_logic_vector) return int777_t is
  variable rv : int777_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint778_t_to_slv(x : uint778_t) return std_logic_vector is
  variable rv : std_logic_vector(777 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint778_t(x : std_logic_vector) return uint778_t is
  variable rv : uint778_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int778_t_to_slv(x : int778_t) return std_logic_vector is
  variable rv : std_logic_vector(777 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int778_t(x : std_logic_vector) return int778_t is
  variable rv : int778_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint779_t_to_slv(x : uint779_t) return std_logic_vector is
  variable rv : std_logic_vector(778 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint779_t(x : std_logic_vector) return uint779_t is
  variable rv : uint779_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int779_t_to_slv(x : int779_t) return std_logic_vector is
  variable rv : std_logic_vector(778 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int779_t(x : std_logic_vector) return int779_t is
  variable rv : int779_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint780_t_to_slv(x : uint780_t) return std_logic_vector is
  variable rv : std_logic_vector(779 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint780_t(x : std_logic_vector) return uint780_t is
  variable rv : uint780_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int780_t_to_slv(x : int780_t) return std_logic_vector is
  variable rv : std_logic_vector(779 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int780_t(x : std_logic_vector) return int780_t is
  variable rv : int780_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint781_t_to_slv(x : uint781_t) return std_logic_vector is
  variable rv : std_logic_vector(780 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint781_t(x : std_logic_vector) return uint781_t is
  variable rv : uint781_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int781_t_to_slv(x : int781_t) return std_logic_vector is
  variable rv : std_logic_vector(780 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int781_t(x : std_logic_vector) return int781_t is
  variable rv : int781_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint782_t_to_slv(x : uint782_t) return std_logic_vector is
  variable rv : std_logic_vector(781 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint782_t(x : std_logic_vector) return uint782_t is
  variable rv : uint782_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int782_t_to_slv(x : int782_t) return std_logic_vector is
  variable rv : std_logic_vector(781 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int782_t(x : std_logic_vector) return int782_t is
  variable rv : int782_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint783_t_to_slv(x : uint783_t) return std_logic_vector is
  variable rv : std_logic_vector(782 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint783_t(x : std_logic_vector) return uint783_t is
  variable rv : uint783_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int783_t_to_slv(x : int783_t) return std_logic_vector is
  variable rv : std_logic_vector(782 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int783_t(x : std_logic_vector) return int783_t is
  variable rv : int783_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint784_t_to_slv(x : uint784_t) return std_logic_vector is
  variable rv : std_logic_vector(783 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint784_t(x : std_logic_vector) return uint784_t is
  variable rv : uint784_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int784_t_to_slv(x : int784_t) return std_logic_vector is
  variable rv : std_logic_vector(783 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int784_t(x : std_logic_vector) return int784_t is
  variable rv : int784_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint785_t_to_slv(x : uint785_t) return std_logic_vector is
  variable rv : std_logic_vector(784 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint785_t(x : std_logic_vector) return uint785_t is
  variable rv : uint785_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int785_t_to_slv(x : int785_t) return std_logic_vector is
  variable rv : std_logic_vector(784 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int785_t(x : std_logic_vector) return int785_t is
  variable rv : int785_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint786_t_to_slv(x : uint786_t) return std_logic_vector is
  variable rv : std_logic_vector(785 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint786_t(x : std_logic_vector) return uint786_t is
  variable rv : uint786_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int786_t_to_slv(x : int786_t) return std_logic_vector is
  variable rv : std_logic_vector(785 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int786_t(x : std_logic_vector) return int786_t is
  variable rv : int786_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint787_t_to_slv(x : uint787_t) return std_logic_vector is
  variable rv : std_logic_vector(786 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint787_t(x : std_logic_vector) return uint787_t is
  variable rv : uint787_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int787_t_to_slv(x : int787_t) return std_logic_vector is
  variable rv : std_logic_vector(786 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int787_t(x : std_logic_vector) return int787_t is
  variable rv : int787_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint788_t_to_slv(x : uint788_t) return std_logic_vector is
  variable rv : std_logic_vector(787 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint788_t(x : std_logic_vector) return uint788_t is
  variable rv : uint788_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int788_t_to_slv(x : int788_t) return std_logic_vector is
  variable rv : std_logic_vector(787 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int788_t(x : std_logic_vector) return int788_t is
  variable rv : int788_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint789_t_to_slv(x : uint789_t) return std_logic_vector is
  variable rv : std_logic_vector(788 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint789_t(x : std_logic_vector) return uint789_t is
  variable rv : uint789_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int789_t_to_slv(x : int789_t) return std_logic_vector is
  variable rv : std_logic_vector(788 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int789_t(x : std_logic_vector) return int789_t is
  variable rv : int789_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint790_t_to_slv(x : uint790_t) return std_logic_vector is
  variable rv : std_logic_vector(789 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint790_t(x : std_logic_vector) return uint790_t is
  variable rv : uint790_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int790_t_to_slv(x : int790_t) return std_logic_vector is
  variable rv : std_logic_vector(789 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int790_t(x : std_logic_vector) return int790_t is
  variable rv : int790_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint791_t_to_slv(x : uint791_t) return std_logic_vector is
  variable rv : std_logic_vector(790 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint791_t(x : std_logic_vector) return uint791_t is
  variable rv : uint791_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int791_t_to_slv(x : int791_t) return std_logic_vector is
  variable rv : std_logic_vector(790 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int791_t(x : std_logic_vector) return int791_t is
  variable rv : int791_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint792_t_to_slv(x : uint792_t) return std_logic_vector is
  variable rv : std_logic_vector(791 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint792_t(x : std_logic_vector) return uint792_t is
  variable rv : uint792_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int792_t_to_slv(x : int792_t) return std_logic_vector is
  variable rv : std_logic_vector(791 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int792_t(x : std_logic_vector) return int792_t is
  variable rv : int792_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint793_t_to_slv(x : uint793_t) return std_logic_vector is
  variable rv : std_logic_vector(792 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint793_t(x : std_logic_vector) return uint793_t is
  variable rv : uint793_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int793_t_to_slv(x : int793_t) return std_logic_vector is
  variable rv : std_logic_vector(792 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int793_t(x : std_logic_vector) return int793_t is
  variable rv : int793_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint794_t_to_slv(x : uint794_t) return std_logic_vector is
  variable rv : std_logic_vector(793 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint794_t(x : std_logic_vector) return uint794_t is
  variable rv : uint794_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int794_t_to_slv(x : int794_t) return std_logic_vector is
  variable rv : std_logic_vector(793 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int794_t(x : std_logic_vector) return int794_t is
  variable rv : int794_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint795_t_to_slv(x : uint795_t) return std_logic_vector is
  variable rv : std_logic_vector(794 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint795_t(x : std_logic_vector) return uint795_t is
  variable rv : uint795_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int795_t_to_slv(x : int795_t) return std_logic_vector is
  variable rv : std_logic_vector(794 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int795_t(x : std_logic_vector) return int795_t is
  variable rv : int795_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint796_t_to_slv(x : uint796_t) return std_logic_vector is
  variable rv : std_logic_vector(795 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint796_t(x : std_logic_vector) return uint796_t is
  variable rv : uint796_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int796_t_to_slv(x : int796_t) return std_logic_vector is
  variable rv : std_logic_vector(795 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int796_t(x : std_logic_vector) return int796_t is
  variable rv : int796_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint797_t_to_slv(x : uint797_t) return std_logic_vector is
  variable rv : std_logic_vector(796 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint797_t(x : std_logic_vector) return uint797_t is
  variable rv : uint797_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int797_t_to_slv(x : int797_t) return std_logic_vector is
  variable rv : std_logic_vector(796 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int797_t(x : std_logic_vector) return int797_t is
  variable rv : int797_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint798_t_to_slv(x : uint798_t) return std_logic_vector is
  variable rv : std_logic_vector(797 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint798_t(x : std_logic_vector) return uint798_t is
  variable rv : uint798_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int798_t_to_slv(x : int798_t) return std_logic_vector is
  variable rv : std_logic_vector(797 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int798_t(x : std_logic_vector) return int798_t is
  variable rv : int798_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint799_t_to_slv(x : uint799_t) return std_logic_vector is
  variable rv : std_logic_vector(798 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint799_t(x : std_logic_vector) return uint799_t is
  variable rv : uint799_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int799_t_to_slv(x : int799_t) return std_logic_vector is
  variable rv : std_logic_vector(798 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int799_t(x : std_logic_vector) return int799_t is
  variable rv : int799_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint800_t_to_slv(x : uint800_t) return std_logic_vector is
  variable rv : std_logic_vector(799 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint800_t(x : std_logic_vector) return uint800_t is
  variable rv : uint800_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int800_t_to_slv(x : int800_t) return std_logic_vector is
  variable rv : std_logic_vector(799 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int800_t(x : std_logic_vector) return int800_t is
  variable rv : int800_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint801_t_to_slv(x : uint801_t) return std_logic_vector is
  variable rv : std_logic_vector(800 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint801_t(x : std_logic_vector) return uint801_t is
  variable rv : uint801_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int801_t_to_slv(x : int801_t) return std_logic_vector is
  variable rv : std_logic_vector(800 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int801_t(x : std_logic_vector) return int801_t is
  variable rv : int801_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint802_t_to_slv(x : uint802_t) return std_logic_vector is
  variable rv : std_logic_vector(801 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint802_t(x : std_logic_vector) return uint802_t is
  variable rv : uint802_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int802_t_to_slv(x : int802_t) return std_logic_vector is
  variable rv : std_logic_vector(801 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int802_t(x : std_logic_vector) return int802_t is
  variable rv : int802_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint803_t_to_slv(x : uint803_t) return std_logic_vector is
  variable rv : std_logic_vector(802 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint803_t(x : std_logic_vector) return uint803_t is
  variable rv : uint803_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int803_t_to_slv(x : int803_t) return std_logic_vector is
  variable rv : std_logic_vector(802 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int803_t(x : std_logic_vector) return int803_t is
  variable rv : int803_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint804_t_to_slv(x : uint804_t) return std_logic_vector is
  variable rv : std_logic_vector(803 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint804_t(x : std_logic_vector) return uint804_t is
  variable rv : uint804_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int804_t_to_slv(x : int804_t) return std_logic_vector is
  variable rv : std_logic_vector(803 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int804_t(x : std_logic_vector) return int804_t is
  variable rv : int804_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint805_t_to_slv(x : uint805_t) return std_logic_vector is
  variable rv : std_logic_vector(804 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint805_t(x : std_logic_vector) return uint805_t is
  variable rv : uint805_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int805_t_to_slv(x : int805_t) return std_logic_vector is
  variable rv : std_logic_vector(804 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int805_t(x : std_logic_vector) return int805_t is
  variable rv : int805_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint806_t_to_slv(x : uint806_t) return std_logic_vector is
  variable rv : std_logic_vector(805 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint806_t(x : std_logic_vector) return uint806_t is
  variable rv : uint806_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int806_t_to_slv(x : int806_t) return std_logic_vector is
  variable rv : std_logic_vector(805 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int806_t(x : std_logic_vector) return int806_t is
  variable rv : int806_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint807_t_to_slv(x : uint807_t) return std_logic_vector is
  variable rv : std_logic_vector(806 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint807_t(x : std_logic_vector) return uint807_t is
  variable rv : uint807_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int807_t_to_slv(x : int807_t) return std_logic_vector is
  variable rv : std_logic_vector(806 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int807_t(x : std_logic_vector) return int807_t is
  variable rv : int807_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint808_t_to_slv(x : uint808_t) return std_logic_vector is
  variable rv : std_logic_vector(807 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint808_t(x : std_logic_vector) return uint808_t is
  variable rv : uint808_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int808_t_to_slv(x : int808_t) return std_logic_vector is
  variable rv : std_logic_vector(807 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int808_t(x : std_logic_vector) return int808_t is
  variable rv : int808_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint809_t_to_slv(x : uint809_t) return std_logic_vector is
  variable rv : std_logic_vector(808 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint809_t(x : std_logic_vector) return uint809_t is
  variable rv : uint809_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int809_t_to_slv(x : int809_t) return std_logic_vector is
  variable rv : std_logic_vector(808 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int809_t(x : std_logic_vector) return int809_t is
  variable rv : int809_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint810_t_to_slv(x : uint810_t) return std_logic_vector is
  variable rv : std_logic_vector(809 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint810_t(x : std_logic_vector) return uint810_t is
  variable rv : uint810_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int810_t_to_slv(x : int810_t) return std_logic_vector is
  variable rv : std_logic_vector(809 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int810_t(x : std_logic_vector) return int810_t is
  variable rv : int810_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint811_t_to_slv(x : uint811_t) return std_logic_vector is
  variable rv : std_logic_vector(810 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint811_t(x : std_logic_vector) return uint811_t is
  variable rv : uint811_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int811_t_to_slv(x : int811_t) return std_logic_vector is
  variable rv : std_logic_vector(810 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int811_t(x : std_logic_vector) return int811_t is
  variable rv : int811_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint812_t_to_slv(x : uint812_t) return std_logic_vector is
  variable rv : std_logic_vector(811 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint812_t(x : std_logic_vector) return uint812_t is
  variable rv : uint812_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int812_t_to_slv(x : int812_t) return std_logic_vector is
  variable rv : std_logic_vector(811 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int812_t(x : std_logic_vector) return int812_t is
  variable rv : int812_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint813_t_to_slv(x : uint813_t) return std_logic_vector is
  variable rv : std_logic_vector(812 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint813_t(x : std_logic_vector) return uint813_t is
  variable rv : uint813_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int813_t_to_slv(x : int813_t) return std_logic_vector is
  variable rv : std_logic_vector(812 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int813_t(x : std_logic_vector) return int813_t is
  variable rv : int813_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint814_t_to_slv(x : uint814_t) return std_logic_vector is
  variable rv : std_logic_vector(813 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint814_t(x : std_logic_vector) return uint814_t is
  variable rv : uint814_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int814_t_to_slv(x : int814_t) return std_logic_vector is
  variable rv : std_logic_vector(813 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int814_t(x : std_logic_vector) return int814_t is
  variable rv : int814_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint815_t_to_slv(x : uint815_t) return std_logic_vector is
  variable rv : std_logic_vector(814 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint815_t(x : std_logic_vector) return uint815_t is
  variable rv : uint815_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int815_t_to_slv(x : int815_t) return std_logic_vector is
  variable rv : std_logic_vector(814 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int815_t(x : std_logic_vector) return int815_t is
  variable rv : int815_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint816_t_to_slv(x : uint816_t) return std_logic_vector is
  variable rv : std_logic_vector(815 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint816_t(x : std_logic_vector) return uint816_t is
  variable rv : uint816_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int816_t_to_slv(x : int816_t) return std_logic_vector is
  variable rv : std_logic_vector(815 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int816_t(x : std_logic_vector) return int816_t is
  variable rv : int816_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint817_t_to_slv(x : uint817_t) return std_logic_vector is
  variable rv : std_logic_vector(816 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint817_t(x : std_logic_vector) return uint817_t is
  variable rv : uint817_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int817_t_to_slv(x : int817_t) return std_logic_vector is
  variable rv : std_logic_vector(816 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int817_t(x : std_logic_vector) return int817_t is
  variable rv : int817_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint818_t_to_slv(x : uint818_t) return std_logic_vector is
  variable rv : std_logic_vector(817 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint818_t(x : std_logic_vector) return uint818_t is
  variable rv : uint818_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int818_t_to_slv(x : int818_t) return std_logic_vector is
  variable rv : std_logic_vector(817 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int818_t(x : std_logic_vector) return int818_t is
  variable rv : int818_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint819_t_to_slv(x : uint819_t) return std_logic_vector is
  variable rv : std_logic_vector(818 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint819_t(x : std_logic_vector) return uint819_t is
  variable rv : uint819_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int819_t_to_slv(x : int819_t) return std_logic_vector is
  variable rv : std_logic_vector(818 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int819_t(x : std_logic_vector) return int819_t is
  variable rv : int819_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint820_t_to_slv(x : uint820_t) return std_logic_vector is
  variable rv : std_logic_vector(819 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint820_t(x : std_logic_vector) return uint820_t is
  variable rv : uint820_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int820_t_to_slv(x : int820_t) return std_logic_vector is
  variable rv : std_logic_vector(819 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int820_t(x : std_logic_vector) return int820_t is
  variable rv : int820_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint821_t_to_slv(x : uint821_t) return std_logic_vector is
  variable rv : std_logic_vector(820 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint821_t(x : std_logic_vector) return uint821_t is
  variable rv : uint821_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int821_t_to_slv(x : int821_t) return std_logic_vector is
  variable rv : std_logic_vector(820 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int821_t(x : std_logic_vector) return int821_t is
  variable rv : int821_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint822_t_to_slv(x : uint822_t) return std_logic_vector is
  variable rv : std_logic_vector(821 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint822_t(x : std_logic_vector) return uint822_t is
  variable rv : uint822_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int822_t_to_slv(x : int822_t) return std_logic_vector is
  variable rv : std_logic_vector(821 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int822_t(x : std_logic_vector) return int822_t is
  variable rv : int822_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint823_t_to_slv(x : uint823_t) return std_logic_vector is
  variable rv : std_logic_vector(822 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint823_t(x : std_logic_vector) return uint823_t is
  variable rv : uint823_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int823_t_to_slv(x : int823_t) return std_logic_vector is
  variable rv : std_logic_vector(822 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int823_t(x : std_logic_vector) return int823_t is
  variable rv : int823_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint824_t_to_slv(x : uint824_t) return std_logic_vector is
  variable rv : std_logic_vector(823 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint824_t(x : std_logic_vector) return uint824_t is
  variable rv : uint824_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int824_t_to_slv(x : int824_t) return std_logic_vector is
  variable rv : std_logic_vector(823 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int824_t(x : std_logic_vector) return int824_t is
  variable rv : int824_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint825_t_to_slv(x : uint825_t) return std_logic_vector is
  variable rv : std_logic_vector(824 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint825_t(x : std_logic_vector) return uint825_t is
  variable rv : uint825_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int825_t_to_slv(x : int825_t) return std_logic_vector is
  variable rv : std_logic_vector(824 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int825_t(x : std_logic_vector) return int825_t is
  variable rv : int825_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint826_t_to_slv(x : uint826_t) return std_logic_vector is
  variable rv : std_logic_vector(825 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint826_t(x : std_logic_vector) return uint826_t is
  variable rv : uint826_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int826_t_to_slv(x : int826_t) return std_logic_vector is
  variable rv : std_logic_vector(825 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int826_t(x : std_logic_vector) return int826_t is
  variable rv : int826_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint827_t_to_slv(x : uint827_t) return std_logic_vector is
  variable rv : std_logic_vector(826 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint827_t(x : std_logic_vector) return uint827_t is
  variable rv : uint827_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int827_t_to_slv(x : int827_t) return std_logic_vector is
  variable rv : std_logic_vector(826 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int827_t(x : std_logic_vector) return int827_t is
  variable rv : int827_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint828_t_to_slv(x : uint828_t) return std_logic_vector is
  variable rv : std_logic_vector(827 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint828_t(x : std_logic_vector) return uint828_t is
  variable rv : uint828_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int828_t_to_slv(x : int828_t) return std_logic_vector is
  variable rv : std_logic_vector(827 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int828_t(x : std_logic_vector) return int828_t is
  variable rv : int828_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint829_t_to_slv(x : uint829_t) return std_logic_vector is
  variable rv : std_logic_vector(828 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint829_t(x : std_logic_vector) return uint829_t is
  variable rv : uint829_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int829_t_to_slv(x : int829_t) return std_logic_vector is
  variable rv : std_logic_vector(828 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int829_t(x : std_logic_vector) return int829_t is
  variable rv : int829_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint830_t_to_slv(x : uint830_t) return std_logic_vector is
  variable rv : std_logic_vector(829 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint830_t(x : std_logic_vector) return uint830_t is
  variable rv : uint830_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int830_t_to_slv(x : int830_t) return std_logic_vector is
  variable rv : std_logic_vector(829 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int830_t(x : std_logic_vector) return int830_t is
  variable rv : int830_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint831_t_to_slv(x : uint831_t) return std_logic_vector is
  variable rv : std_logic_vector(830 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint831_t(x : std_logic_vector) return uint831_t is
  variable rv : uint831_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int831_t_to_slv(x : int831_t) return std_logic_vector is
  variable rv : std_logic_vector(830 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int831_t(x : std_logic_vector) return int831_t is
  variable rv : int831_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint832_t_to_slv(x : uint832_t) return std_logic_vector is
  variable rv : std_logic_vector(831 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint832_t(x : std_logic_vector) return uint832_t is
  variable rv : uint832_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int832_t_to_slv(x : int832_t) return std_logic_vector is
  variable rv : std_logic_vector(831 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int832_t(x : std_logic_vector) return int832_t is
  variable rv : int832_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint833_t_to_slv(x : uint833_t) return std_logic_vector is
  variable rv : std_logic_vector(832 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint833_t(x : std_logic_vector) return uint833_t is
  variable rv : uint833_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int833_t_to_slv(x : int833_t) return std_logic_vector is
  variable rv : std_logic_vector(832 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int833_t(x : std_logic_vector) return int833_t is
  variable rv : int833_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint834_t_to_slv(x : uint834_t) return std_logic_vector is
  variable rv : std_logic_vector(833 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint834_t(x : std_logic_vector) return uint834_t is
  variable rv : uint834_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int834_t_to_slv(x : int834_t) return std_logic_vector is
  variable rv : std_logic_vector(833 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int834_t(x : std_logic_vector) return int834_t is
  variable rv : int834_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint835_t_to_slv(x : uint835_t) return std_logic_vector is
  variable rv : std_logic_vector(834 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint835_t(x : std_logic_vector) return uint835_t is
  variable rv : uint835_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int835_t_to_slv(x : int835_t) return std_logic_vector is
  variable rv : std_logic_vector(834 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int835_t(x : std_logic_vector) return int835_t is
  variable rv : int835_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint836_t_to_slv(x : uint836_t) return std_logic_vector is
  variable rv : std_logic_vector(835 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint836_t(x : std_logic_vector) return uint836_t is
  variable rv : uint836_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int836_t_to_slv(x : int836_t) return std_logic_vector is
  variable rv : std_logic_vector(835 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int836_t(x : std_logic_vector) return int836_t is
  variable rv : int836_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint837_t_to_slv(x : uint837_t) return std_logic_vector is
  variable rv : std_logic_vector(836 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint837_t(x : std_logic_vector) return uint837_t is
  variable rv : uint837_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int837_t_to_slv(x : int837_t) return std_logic_vector is
  variable rv : std_logic_vector(836 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int837_t(x : std_logic_vector) return int837_t is
  variable rv : int837_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint838_t_to_slv(x : uint838_t) return std_logic_vector is
  variable rv : std_logic_vector(837 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint838_t(x : std_logic_vector) return uint838_t is
  variable rv : uint838_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int838_t_to_slv(x : int838_t) return std_logic_vector is
  variable rv : std_logic_vector(837 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int838_t(x : std_logic_vector) return int838_t is
  variable rv : int838_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint839_t_to_slv(x : uint839_t) return std_logic_vector is
  variable rv : std_logic_vector(838 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint839_t(x : std_logic_vector) return uint839_t is
  variable rv : uint839_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int839_t_to_slv(x : int839_t) return std_logic_vector is
  variable rv : std_logic_vector(838 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int839_t(x : std_logic_vector) return int839_t is
  variable rv : int839_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint840_t_to_slv(x : uint840_t) return std_logic_vector is
  variable rv : std_logic_vector(839 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint840_t(x : std_logic_vector) return uint840_t is
  variable rv : uint840_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int840_t_to_slv(x : int840_t) return std_logic_vector is
  variable rv : std_logic_vector(839 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int840_t(x : std_logic_vector) return int840_t is
  variable rv : int840_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint841_t_to_slv(x : uint841_t) return std_logic_vector is
  variable rv : std_logic_vector(840 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint841_t(x : std_logic_vector) return uint841_t is
  variable rv : uint841_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int841_t_to_slv(x : int841_t) return std_logic_vector is
  variable rv : std_logic_vector(840 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int841_t(x : std_logic_vector) return int841_t is
  variable rv : int841_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint842_t_to_slv(x : uint842_t) return std_logic_vector is
  variable rv : std_logic_vector(841 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint842_t(x : std_logic_vector) return uint842_t is
  variable rv : uint842_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int842_t_to_slv(x : int842_t) return std_logic_vector is
  variable rv : std_logic_vector(841 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int842_t(x : std_logic_vector) return int842_t is
  variable rv : int842_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint843_t_to_slv(x : uint843_t) return std_logic_vector is
  variable rv : std_logic_vector(842 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint843_t(x : std_logic_vector) return uint843_t is
  variable rv : uint843_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int843_t_to_slv(x : int843_t) return std_logic_vector is
  variable rv : std_logic_vector(842 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int843_t(x : std_logic_vector) return int843_t is
  variable rv : int843_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint844_t_to_slv(x : uint844_t) return std_logic_vector is
  variable rv : std_logic_vector(843 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint844_t(x : std_logic_vector) return uint844_t is
  variable rv : uint844_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int844_t_to_slv(x : int844_t) return std_logic_vector is
  variable rv : std_logic_vector(843 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int844_t(x : std_logic_vector) return int844_t is
  variable rv : int844_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint845_t_to_slv(x : uint845_t) return std_logic_vector is
  variable rv : std_logic_vector(844 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint845_t(x : std_logic_vector) return uint845_t is
  variable rv : uint845_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int845_t_to_slv(x : int845_t) return std_logic_vector is
  variable rv : std_logic_vector(844 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int845_t(x : std_logic_vector) return int845_t is
  variable rv : int845_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint846_t_to_slv(x : uint846_t) return std_logic_vector is
  variable rv : std_logic_vector(845 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint846_t(x : std_logic_vector) return uint846_t is
  variable rv : uint846_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int846_t_to_slv(x : int846_t) return std_logic_vector is
  variable rv : std_logic_vector(845 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int846_t(x : std_logic_vector) return int846_t is
  variable rv : int846_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint847_t_to_slv(x : uint847_t) return std_logic_vector is
  variable rv : std_logic_vector(846 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint847_t(x : std_logic_vector) return uint847_t is
  variable rv : uint847_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int847_t_to_slv(x : int847_t) return std_logic_vector is
  variable rv : std_logic_vector(846 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int847_t(x : std_logic_vector) return int847_t is
  variable rv : int847_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint848_t_to_slv(x : uint848_t) return std_logic_vector is
  variable rv : std_logic_vector(847 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint848_t(x : std_logic_vector) return uint848_t is
  variable rv : uint848_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int848_t_to_slv(x : int848_t) return std_logic_vector is
  variable rv : std_logic_vector(847 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int848_t(x : std_logic_vector) return int848_t is
  variable rv : int848_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint849_t_to_slv(x : uint849_t) return std_logic_vector is
  variable rv : std_logic_vector(848 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint849_t(x : std_logic_vector) return uint849_t is
  variable rv : uint849_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int849_t_to_slv(x : int849_t) return std_logic_vector is
  variable rv : std_logic_vector(848 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int849_t(x : std_logic_vector) return int849_t is
  variable rv : int849_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint850_t_to_slv(x : uint850_t) return std_logic_vector is
  variable rv : std_logic_vector(849 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint850_t(x : std_logic_vector) return uint850_t is
  variable rv : uint850_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int850_t_to_slv(x : int850_t) return std_logic_vector is
  variable rv : std_logic_vector(849 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int850_t(x : std_logic_vector) return int850_t is
  variable rv : int850_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint851_t_to_slv(x : uint851_t) return std_logic_vector is
  variable rv : std_logic_vector(850 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint851_t(x : std_logic_vector) return uint851_t is
  variable rv : uint851_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int851_t_to_slv(x : int851_t) return std_logic_vector is
  variable rv : std_logic_vector(850 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int851_t(x : std_logic_vector) return int851_t is
  variable rv : int851_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint852_t_to_slv(x : uint852_t) return std_logic_vector is
  variable rv : std_logic_vector(851 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint852_t(x : std_logic_vector) return uint852_t is
  variable rv : uint852_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int852_t_to_slv(x : int852_t) return std_logic_vector is
  variable rv : std_logic_vector(851 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int852_t(x : std_logic_vector) return int852_t is
  variable rv : int852_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint853_t_to_slv(x : uint853_t) return std_logic_vector is
  variable rv : std_logic_vector(852 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint853_t(x : std_logic_vector) return uint853_t is
  variable rv : uint853_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int853_t_to_slv(x : int853_t) return std_logic_vector is
  variable rv : std_logic_vector(852 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int853_t(x : std_logic_vector) return int853_t is
  variable rv : int853_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint854_t_to_slv(x : uint854_t) return std_logic_vector is
  variable rv : std_logic_vector(853 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint854_t(x : std_logic_vector) return uint854_t is
  variable rv : uint854_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int854_t_to_slv(x : int854_t) return std_logic_vector is
  variable rv : std_logic_vector(853 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int854_t(x : std_logic_vector) return int854_t is
  variable rv : int854_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint855_t_to_slv(x : uint855_t) return std_logic_vector is
  variable rv : std_logic_vector(854 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint855_t(x : std_logic_vector) return uint855_t is
  variable rv : uint855_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int855_t_to_slv(x : int855_t) return std_logic_vector is
  variable rv : std_logic_vector(854 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int855_t(x : std_logic_vector) return int855_t is
  variable rv : int855_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint856_t_to_slv(x : uint856_t) return std_logic_vector is
  variable rv : std_logic_vector(855 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint856_t(x : std_logic_vector) return uint856_t is
  variable rv : uint856_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int856_t_to_slv(x : int856_t) return std_logic_vector is
  variable rv : std_logic_vector(855 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int856_t(x : std_logic_vector) return int856_t is
  variable rv : int856_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint857_t_to_slv(x : uint857_t) return std_logic_vector is
  variable rv : std_logic_vector(856 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint857_t(x : std_logic_vector) return uint857_t is
  variable rv : uint857_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int857_t_to_slv(x : int857_t) return std_logic_vector is
  variable rv : std_logic_vector(856 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int857_t(x : std_logic_vector) return int857_t is
  variable rv : int857_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint858_t_to_slv(x : uint858_t) return std_logic_vector is
  variable rv : std_logic_vector(857 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint858_t(x : std_logic_vector) return uint858_t is
  variable rv : uint858_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int858_t_to_slv(x : int858_t) return std_logic_vector is
  variable rv : std_logic_vector(857 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int858_t(x : std_logic_vector) return int858_t is
  variable rv : int858_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint859_t_to_slv(x : uint859_t) return std_logic_vector is
  variable rv : std_logic_vector(858 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint859_t(x : std_logic_vector) return uint859_t is
  variable rv : uint859_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int859_t_to_slv(x : int859_t) return std_logic_vector is
  variable rv : std_logic_vector(858 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int859_t(x : std_logic_vector) return int859_t is
  variable rv : int859_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint860_t_to_slv(x : uint860_t) return std_logic_vector is
  variable rv : std_logic_vector(859 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint860_t(x : std_logic_vector) return uint860_t is
  variable rv : uint860_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int860_t_to_slv(x : int860_t) return std_logic_vector is
  variable rv : std_logic_vector(859 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int860_t(x : std_logic_vector) return int860_t is
  variable rv : int860_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint861_t_to_slv(x : uint861_t) return std_logic_vector is
  variable rv : std_logic_vector(860 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint861_t(x : std_logic_vector) return uint861_t is
  variable rv : uint861_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int861_t_to_slv(x : int861_t) return std_logic_vector is
  variable rv : std_logic_vector(860 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int861_t(x : std_logic_vector) return int861_t is
  variable rv : int861_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint862_t_to_slv(x : uint862_t) return std_logic_vector is
  variable rv : std_logic_vector(861 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint862_t(x : std_logic_vector) return uint862_t is
  variable rv : uint862_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int862_t_to_slv(x : int862_t) return std_logic_vector is
  variable rv : std_logic_vector(861 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int862_t(x : std_logic_vector) return int862_t is
  variable rv : int862_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint863_t_to_slv(x : uint863_t) return std_logic_vector is
  variable rv : std_logic_vector(862 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint863_t(x : std_logic_vector) return uint863_t is
  variable rv : uint863_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int863_t_to_slv(x : int863_t) return std_logic_vector is
  variable rv : std_logic_vector(862 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int863_t(x : std_logic_vector) return int863_t is
  variable rv : int863_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint864_t_to_slv(x : uint864_t) return std_logic_vector is
  variable rv : std_logic_vector(863 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint864_t(x : std_logic_vector) return uint864_t is
  variable rv : uint864_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int864_t_to_slv(x : int864_t) return std_logic_vector is
  variable rv : std_logic_vector(863 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int864_t(x : std_logic_vector) return int864_t is
  variable rv : int864_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint865_t_to_slv(x : uint865_t) return std_logic_vector is
  variable rv : std_logic_vector(864 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint865_t(x : std_logic_vector) return uint865_t is
  variable rv : uint865_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int865_t_to_slv(x : int865_t) return std_logic_vector is
  variable rv : std_logic_vector(864 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int865_t(x : std_logic_vector) return int865_t is
  variable rv : int865_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint866_t_to_slv(x : uint866_t) return std_logic_vector is
  variable rv : std_logic_vector(865 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint866_t(x : std_logic_vector) return uint866_t is
  variable rv : uint866_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int866_t_to_slv(x : int866_t) return std_logic_vector is
  variable rv : std_logic_vector(865 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int866_t(x : std_logic_vector) return int866_t is
  variable rv : int866_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint867_t_to_slv(x : uint867_t) return std_logic_vector is
  variable rv : std_logic_vector(866 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint867_t(x : std_logic_vector) return uint867_t is
  variable rv : uint867_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int867_t_to_slv(x : int867_t) return std_logic_vector is
  variable rv : std_logic_vector(866 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int867_t(x : std_logic_vector) return int867_t is
  variable rv : int867_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint868_t_to_slv(x : uint868_t) return std_logic_vector is
  variable rv : std_logic_vector(867 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint868_t(x : std_logic_vector) return uint868_t is
  variable rv : uint868_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int868_t_to_slv(x : int868_t) return std_logic_vector is
  variable rv : std_logic_vector(867 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int868_t(x : std_logic_vector) return int868_t is
  variable rv : int868_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint869_t_to_slv(x : uint869_t) return std_logic_vector is
  variable rv : std_logic_vector(868 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint869_t(x : std_logic_vector) return uint869_t is
  variable rv : uint869_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int869_t_to_slv(x : int869_t) return std_logic_vector is
  variable rv : std_logic_vector(868 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int869_t(x : std_logic_vector) return int869_t is
  variable rv : int869_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint870_t_to_slv(x : uint870_t) return std_logic_vector is
  variable rv : std_logic_vector(869 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint870_t(x : std_logic_vector) return uint870_t is
  variable rv : uint870_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int870_t_to_slv(x : int870_t) return std_logic_vector is
  variable rv : std_logic_vector(869 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int870_t(x : std_logic_vector) return int870_t is
  variable rv : int870_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint871_t_to_slv(x : uint871_t) return std_logic_vector is
  variable rv : std_logic_vector(870 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint871_t(x : std_logic_vector) return uint871_t is
  variable rv : uint871_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int871_t_to_slv(x : int871_t) return std_logic_vector is
  variable rv : std_logic_vector(870 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int871_t(x : std_logic_vector) return int871_t is
  variable rv : int871_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint872_t_to_slv(x : uint872_t) return std_logic_vector is
  variable rv : std_logic_vector(871 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint872_t(x : std_logic_vector) return uint872_t is
  variable rv : uint872_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int872_t_to_slv(x : int872_t) return std_logic_vector is
  variable rv : std_logic_vector(871 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int872_t(x : std_logic_vector) return int872_t is
  variable rv : int872_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint873_t_to_slv(x : uint873_t) return std_logic_vector is
  variable rv : std_logic_vector(872 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint873_t(x : std_logic_vector) return uint873_t is
  variable rv : uint873_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int873_t_to_slv(x : int873_t) return std_logic_vector is
  variable rv : std_logic_vector(872 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int873_t(x : std_logic_vector) return int873_t is
  variable rv : int873_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint874_t_to_slv(x : uint874_t) return std_logic_vector is
  variable rv : std_logic_vector(873 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint874_t(x : std_logic_vector) return uint874_t is
  variable rv : uint874_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int874_t_to_slv(x : int874_t) return std_logic_vector is
  variable rv : std_logic_vector(873 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int874_t(x : std_logic_vector) return int874_t is
  variable rv : int874_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint875_t_to_slv(x : uint875_t) return std_logic_vector is
  variable rv : std_logic_vector(874 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint875_t(x : std_logic_vector) return uint875_t is
  variable rv : uint875_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int875_t_to_slv(x : int875_t) return std_logic_vector is
  variable rv : std_logic_vector(874 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int875_t(x : std_logic_vector) return int875_t is
  variable rv : int875_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint876_t_to_slv(x : uint876_t) return std_logic_vector is
  variable rv : std_logic_vector(875 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint876_t(x : std_logic_vector) return uint876_t is
  variable rv : uint876_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int876_t_to_slv(x : int876_t) return std_logic_vector is
  variable rv : std_logic_vector(875 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int876_t(x : std_logic_vector) return int876_t is
  variable rv : int876_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint877_t_to_slv(x : uint877_t) return std_logic_vector is
  variable rv : std_logic_vector(876 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint877_t(x : std_logic_vector) return uint877_t is
  variable rv : uint877_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int877_t_to_slv(x : int877_t) return std_logic_vector is
  variable rv : std_logic_vector(876 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int877_t(x : std_logic_vector) return int877_t is
  variable rv : int877_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint878_t_to_slv(x : uint878_t) return std_logic_vector is
  variable rv : std_logic_vector(877 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint878_t(x : std_logic_vector) return uint878_t is
  variable rv : uint878_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int878_t_to_slv(x : int878_t) return std_logic_vector is
  variable rv : std_logic_vector(877 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int878_t(x : std_logic_vector) return int878_t is
  variable rv : int878_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint879_t_to_slv(x : uint879_t) return std_logic_vector is
  variable rv : std_logic_vector(878 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint879_t(x : std_logic_vector) return uint879_t is
  variable rv : uint879_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int879_t_to_slv(x : int879_t) return std_logic_vector is
  variable rv : std_logic_vector(878 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int879_t(x : std_logic_vector) return int879_t is
  variable rv : int879_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint880_t_to_slv(x : uint880_t) return std_logic_vector is
  variable rv : std_logic_vector(879 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint880_t(x : std_logic_vector) return uint880_t is
  variable rv : uint880_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int880_t_to_slv(x : int880_t) return std_logic_vector is
  variable rv : std_logic_vector(879 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int880_t(x : std_logic_vector) return int880_t is
  variable rv : int880_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint881_t_to_slv(x : uint881_t) return std_logic_vector is
  variable rv : std_logic_vector(880 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint881_t(x : std_logic_vector) return uint881_t is
  variable rv : uint881_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int881_t_to_slv(x : int881_t) return std_logic_vector is
  variable rv : std_logic_vector(880 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int881_t(x : std_logic_vector) return int881_t is
  variable rv : int881_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint882_t_to_slv(x : uint882_t) return std_logic_vector is
  variable rv : std_logic_vector(881 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint882_t(x : std_logic_vector) return uint882_t is
  variable rv : uint882_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int882_t_to_slv(x : int882_t) return std_logic_vector is
  variable rv : std_logic_vector(881 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int882_t(x : std_logic_vector) return int882_t is
  variable rv : int882_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint883_t_to_slv(x : uint883_t) return std_logic_vector is
  variable rv : std_logic_vector(882 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint883_t(x : std_logic_vector) return uint883_t is
  variable rv : uint883_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int883_t_to_slv(x : int883_t) return std_logic_vector is
  variable rv : std_logic_vector(882 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int883_t(x : std_logic_vector) return int883_t is
  variable rv : int883_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint884_t_to_slv(x : uint884_t) return std_logic_vector is
  variable rv : std_logic_vector(883 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint884_t(x : std_logic_vector) return uint884_t is
  variable rv : uint884_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int884_t_to_slv(x : int884_t) return std_logic_vector is
  variable rv : std_logic_vector(883 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int884_t(x : std_logic_vector) return int884_t is
  variable rv : int884_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint885_t_to_slv(x : uint885_t) return std_logic_vector is
  variable rv : std_logic_vector(884 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint885_t(x : std_logic_vector) return uint885_t is
  variable rv : uint885_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int885_t_to_slv(x : int885_t) return std_logic_vector is
  variable rv : std_logic_vector(884 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int885_t(x : std_logic_vector) return int885_t is
  variable rv : int885_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint886_t_to_slv(x : uint886_t) return std_logic_vector is
  variable rv : std_logic_vector(885 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint886_t(x : std_logic_vector) return uint886_t is
  variable rv : uint886_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int886_t_to_slv(x : int886_t) return std_logic_vector is
  variable rv : std_logic_vector(885 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int886_t(x : std_logic_vector) return int886_t is
  variable rv : int886_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint887_t_to_slv(x : uint887_t) return std_logic_vector is
  variable rv : std_logic_vector(886 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint887_t(x : std_logic_vector) return uint887_t is
  variable rv : uint887_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int887_t_to_slv(x : int887_t) return std_logic_vector is
  variable rv : std_logic_vector(886 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int887_t(x : std_logic_vector) return int887_t is
  variable rv : int887_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint888_t_to_slv(x : uint888_t) return std_logic_vector is
  variable rv : std_logic_vector(887 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint888_t(x : std_logic_vector) return uint888_t is
  variable rv : uint888_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int888_t_to_slv(x : int888_t) return std_logic_vector is
  variable rv : std_logic_vector(887 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int888_t(x : std_logic_vector) return int888_t is
  variable rv : int888_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint889_t_to_slv(x : uint889_t) return std_logic_vector is
  variable rv : std_logic_vector(888 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint889_t(x : std_logic_vector) return uint889_t is
  variable rv : uint889_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int889_t_to_slv(x : int889_t) return std_logic_vector is
  variable rv : std_logic_vector(888 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int889_t(x : std_logic_vector) return int889_t is
  variable rv : int889_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint890_t_to_slv(x : uint890_t) return std_logic_vector is
  variable rv : std_logic_vector(889 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint890_t(x : std_logic_vector) return uint890_t is
  variable rv : uint890_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int890_t_to_slv(x : int890_t) return std_logic_vector is
  variable rv : std_logic_vector(889 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int890_t(x : std_logic_vector) return int890_t is
  variable rv : int890_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint891_t_to_slv(x : uint891_t) return std_logic_vector is
  variable rv : std_logic_vector(890 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint891_t(x : std_logic_vector) return uint891_t is
  variable rv : uint891_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int891_t_to_slv(x : int891_t) return std_logic_vector is
  variable rv : std_logic_vector(890 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int891_t(x : std_logic_vector) return int891_t is
  variable rv : int891_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint892_t_to_slv(x : uint892_t) return std_logic_vector is
  variable rv : std_logic_vector(891 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint892_t(x : std_logic_vector) return uint892_t is
  variable rv : uint892_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int892_t_to_slv(x : int892_t) return std_logic_vector is
  variable rv : std_logic_vector(891 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int892_t(x : std_logic_vector) return int892_t is
  variable rv : int892_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint893_t_to_slv(x : uint893_t) return std_logic_vector is
  variable rv : std_logic_vector(892 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint893_t(x : std_logic_vector) return uint893_t is
  variable rv : uint893_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int893_t_to_slv(x : int893_t) return std_logic_vector is
  variable rv : std_logic_vector(892 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int893_t(x : std_logic_vector) return int893_t is
  variable rv : int893_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint894_t_to_slv(x : uint894_t) return std_logic_vector is
  variable rv : std_logic_vector(893 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint894_t(x : std_logic_vector) return uint894_t is
  variable rv : uint894_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int894_t_to_slv(x : int894_t) return std_logic_vector is
  variable rv : std_logic_vector(893 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int894_t(x : std_logic_vector) return int894_t is
  variable rv : int894_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint895_t_to_slv(x : uint895_t) return std_logic_vector is
  variable rv : std_logic_vector(894 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint895_t(x : std_logic_vector) return uint895_t is
  variable rv : uint895_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int895_t_to_slv(x : int895_t) return std_logic_vector is
  variable rv : std_logic_vector(894 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int895_t(x : std_logic_vector) return int895_t is
  variable rv : int895_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint896_t_to_slv(x : uint896_t) return std_logic_vector is
  variable rv : std_logic_vector(895 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint896_t(x : std_logic_vector) return uint896_t is
  variable rv : uint896_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int896_t_to_slv(x : int896_t) return std_logic_vector is
  variable rv : std_logic_vector(895 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int896_t(x : std_logic_vector) return int896_t is
  variable rv : int896_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint897_t_to_slv(x : uint897_t) return std_logic_vector is
  variable rv : std_logic_vector(896 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint897_t(x : std_logic_vector) return uint897_t is
  variable rv : uint897_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int897_t_to_slv(x : int897_t) return std_logic_vector is
  variable rv : std_logic_vector(896 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int897_t(x : std_logic_vector) return int897_t is
  variable rv : int897_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint898_t_to_slv(x : uint898_t) return std_logic_vector is
  variable rv : std_logic_vector(897 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint898_t(x : std_logic_vector) return uint898_t is
  variable rv : uint898_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int898_t_to_slv(x : int898_t) return std_logic_vector is
  variable rv : std_logic_vector(897 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int898_t(x : std_logic_vector) return int898_t is
  variable rv : int898_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint899_t_to_slv(x : uint899_t) return std_logic_vector is
  variable rv : std_logic_vector(898 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint899_t(x : std_logic_vector) return uint899_t is
  variable rv : uint899_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int899_t_to_slv(x : int899_t) return std_logic_vector is
  variable rv : std_logic_vector(898 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int899_t(x : std_logic_vector) return int899_t is
  variable rv : int899_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint900_t_to_slv(x : uint900_t) return std_logic_vector is
  variable rv : std_logic_vector(899 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint900_t(x : std_logic_vector) return uint900_t is
  variable rv : uint900_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int900_t_to_slv(x : int900_t) return std_logic_vector is
  variable rv : std_logic_vector(899 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int900_t(x : std_logic_vector) return int900_t is
  variable rv : int900_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint901_t_to_slv(x : uint901_t) return std_logic_vector is
  variable rv : std_logic_vector(900 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint901_t(x : std_logic_vector) return uint901_t is
  variable rv : uint901_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int901_t_to_slv(x : int901_t) return std_logic_vector is
  variable rv : std_logic_vector(900 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int901_t(x : std_logic_vector) return int901_t is
  variable rv : int901_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint902_t_to_slv(x : uint902_t) return std_logic_vector is
  variable rv : std_logic_vector(901 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint902_t(x : std_logic_vector) return uint902_t is
  variable rv : uint902_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int902_t_to_slv(x : int902_t) return std_logic_vector is
  variable rv : std_logic_vector(901 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int902_t(x : std_logic_vector) return int902_t is
  variable rv : int902_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint903_t_to_slv(x : uint903_t) return std_logic_vector is
  variable rv : std_logic_vector(902 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint903_t(x : std_logic_vector) return uint903_t is
  variable rv : uint903_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int903_t_to_slv(x : int903_t) return std_logic_vector is
  variable rv : std_logic_vector(902 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int903_t(x : std_logic_vector) return int903_t is
  variable rv : int903_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint904_t_to_slv(x : uint904_t) return std_logic_vector is
  variable rv : std_logic_vector(903 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint904_t(x : std_logic_vector) return uint904_t is
  variable rv : uint904_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int904_t_to_slv(x : int904_t) return std_logic_vector is
  variable rv : std_logic_vector(903 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int904_t(x : std_logic_vector) return int904_t is
  variable rv : int904_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint905_t_to_slv(x : uint905_t) return std_logic_vector is
  variable rv : std_logic_vector(904 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint905_t(x : std_logic_vector) return uint905_t is
  variable rv : uint905_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int905_t_to_slv(x : int905_t) return std_logic_vector is
  variable rv : std_logic_vector(904 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int905_t(x : std_logic_vector) return int905_t is
  variable rv : int905_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint906_t_to_slv(x : uint906_t) return std_logic_vector is
  variable rv : std_logic_vector(905 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint906_t(x : std_logic_vector) return uint906_t is
  variable rv : uint906_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int906_t_to_slv(x : int906_t) return std_logic_vector is
  variable rv : std_logic_vector(905 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int906_t(x : std_logic_vector) return int906_t is
  variable rv : int906_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint907_t_to_slv(x : uint907_t) return std_logic_vector is
  variable rv : std_logic_vector(906 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint907_t(x : std_logic_vector) return uint907_t is
  variable rv : uint907_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int907_t_to_slv(x : int907_t) return std_logic_vector is
  variable rv : std_logic_vector(906 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int907_t(x : std_logic_vector) return int907_t is
  variable rv : int907_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint908_t_to_slv(x : uint908_t) return std_logic_vector is
  variable rv : std_logic_vector(907 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint908_t(x : std_logic_vector) return uint908_t is
  variable rv : uint908_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int908_t_to_slv(x : int908_t) return std_logic_vector is
  variable rv : std_logic_vector(907 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int908_t(x : std_logic_vector) return int908_t is
  variable rv : int908_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint909_t_to_slv(x : uint909_t) return std_logic_vector is
  variable rv : std_logic_vector(908 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint909_t(x : std_logic_vector) return uint909_t is
  variable rv : uint909_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int909_t_to_slv(x : int909_t) return std_logic_vector is
  variable rv : std_logic_vector(908 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int909_t(x : std_logic_vector) return int909_t is
  variable rv : int909_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint910_t_to_slv(x : uint910_t) return std_logic_vector is
  variable rv : std_logic_vector(909 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint910_t(x : std_logic_vector) return uint910_t is
  variable rv : uint910_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int910_t_to_slv(x : int910_t) return std_logic_vector is
  variable rv : std_logic_vector(909 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int910_t(x : std_logic_vector) return int910_t is
  variable rv : int910_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint911_t_to_slv(x : uint911_t) return std_logic_vector is
  variable rv : std_logic_vector(910 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint911_t(x : std_logic_vector) return uint911_t is
  variable rv : uint911_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int911_t_to_slv(x : int911_t) return std_logic_vector is
  variable rv : std_logic_vector(910 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int911_t(x : std_logic_vector) return int911_t is
  variable rv : int911_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint912_t_to_slv(x : uint912_t) return std_logic_vector is
  variable rv : std_logic_vector(911 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint912_t(x : std_logic_vector) return uint912_t is
  variable rv : uint912_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int912_t_to_slv(x : int912_t) return std_logic_vector is
  variable rv : std_logic_vector(911 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int912_t(x : std_logic_vector) return int912_t is
  variable rv : int912_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint913_t_to_slv(x : uint913_t) return std_logic_vector is
  variable rv : std_logic_vector(912 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint913_t(x : std_logic_vector) return uint913_t is
  variable rv : uint913_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int913_t_to_slv(x : int913_t) return std_logic_vector is
  variable rv : std_logic_vector(912 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int913_t(x : std_logic_vector) return int913_t is
  variable rv : int913_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint914_t_to_slv(x : uint914_t) return std_logic_vector is
  variable rv : std_logic_vector(913 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint914_t(x : std_logic_vector) return uint914_t is
  variable rv : uint914_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int914_t_to_slv(x : int914_t) return std_logic_vector is
  variable rv : std_logic_vector(913 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int914_t(x : std_logic_vector) return int914_t is
  variable rv : int914_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint915_t_to_slv(x : uint915_t) return std_logic_vector is
  variable rv : std_logic_vector(914 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint915_t(x : std_logic_vector) return uint915_t is
  variable rv : uint915_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int915_t_to_slv(x : int915_t) return std_logic_vector is
  variable rv : std_logic_vector(914 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int915_t(x : std_logic_vector) return int915_t is
  variable rv : int915_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint916_t_to_slv(x : uint916_t) return std_logic_vector is
  variable rv : std_logic_vector(915 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint916_t(x : std_logic_vector) return uint916_t is
  variable rv : uint916_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int916_t_to_slv(x : int916_t) return std_logic_vector is
  variable rv : std_logic_vector(915 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int916_t(x : std_logic_vector) return int916_t is
  variable rv : int916_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint917_t_to_slv(x : uint917_t) return std_logic_vector is
  variable rv : std_logic_vector(916 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint917_t(x : std_logic_vector) return uint917_t is
  variable rv : uint917_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int917_t_to_slv(x : int917_t) return std_logic_vector is
  variable rv : std_logic_vector(916 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int917_t(x : std_logic_vector) return int917_t is
  variable rv : int917_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint918_t_to_slv(x : uint918_t) return std_logic_vector is
  variable rv : std_logic_vector(917 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint918_t(x : std_logic_vector) return uint918_t is
  variable rv : uint918_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int918_t_to_slv(x : int918_t) return std_logic_vector is
  variable rv : std_logic_vector(917 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int918_t(x : std_logic_vector) return int918_t is
  variable rv : int918_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint919_t_to_slv(x : uint919_t) return std_logic_vector is
  variable rv : std_logic_vector(918 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint919_t(x : std_logic_vector) return uint919_t is
  variable rv : uint919_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int919_t_to_slv(x : int919_t) return std_logic_vector is
  variable rv : std_logic_vector(918 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int919_t(x : std_logic_vector) return int919_t is
  variable rv : int919_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint920_t_to_slv(x : uint920_t) return std_logic_vector is
  variable rv : std_logic_vector(919 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint920_t(x : std_logic_vector) return uint920_t is
  variable rv : uint920_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int920_t_to_slv(x : int920_t) return std_logic_vector is
  variable rv : std_logic_vector(919 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int920_t(x : std_logic_vector) return int920_t is
  variable rv : int920_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint921_t_to_slv(x : uint921_t) return std_logic_vector is
  variable rv : std_logic_vector(920 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint921_t(x : std_logic_vector) return uint921_t is
  variable rv : uint921_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int921_t_to_slv(x : int921_t) return std_logic_vector is
  variable rv : std_logic_vector(920 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int921_t(x : std_logic_vector) return int921_t is
  variable rv : int921_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint922_t_to_slv(x : uint922_t) return std_logic_vector is
  variable rv : std_logic_vector(921 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint922_t(x : std_logic_vector) return uint922_t is
  variable rv : uint922_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int922_t_to_slv(x : int922_t) return std_logic_vector is
  variable rv : std_logic_vector(921 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int922_t(x : std_logic_vector) return int922_t is
  variable rv : int922_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint923_t_to_slv(x : uint923_t) return std_logic_vector is
  variable rv : std_logic_vector(922 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint923_t(x : std_logic_vector) return uint923_t is
  variable rv : uint923_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int923_t_to_slv(x : int923_t) return std_logic_vector is
  variable rv : std_logic_vector(922 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int923_t(x : std_logic_vector) return int923_t is
  variable rv : int923_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint924_t_to_slv(x : uint924_t) return std_logic_vector is
  variable rv : std_logic_vector(923 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint924_t(x : std_logic_vector) return uint924_t is
  variable rv : uint924_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int924_t_to_slv(x : int924_t) return std_logic_vector is
  variable rv : std_logic_vector(923 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int924_t(x : std_logic_vector) return int924_t is
  variable rv : int924_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint925_t_to_slv(x : uint925_t) return std_logic_vector is
  variable rv : std_logic_vector(924 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint925_t(x : std_logic_vector) return uint925_t is
  variable rv : uint925_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int925_t_to_slv(x : int925_t) return std_logic_vector is
  variable rv : std_logic_vector(924 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int925_t(x : std_logic_vector) return int925_t is
  variable rv : int925_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint926_t_to_slv(x : uint926_t) return std_logic_vector is
  variable rv : std_logic_vector(925 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint926_t(x : std_logic_vector) return uint926_t is
  variable rv : uint926_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int926_t_to_slv(x : int926_t) return std_logic_vector is
  variable rv : std_logic_vector(925 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int926_t(x : std_logic_vector) return int926_t is
  variable rv : int926_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint927_t_to_slv(x : uint927_t) return std_logic_vector is
  variable rv : std_logic_vector(926 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint927_t(x : std_logic_vector) return uint927_t is
  variable rv : uint927_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int927_t_to_slv(x : int927_t) return std_logic_vector is
  variable rv : std_logic_vector(926 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int927_t(x : std_logic_vector) return int927_t is
  variable rv : int927_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint928_t_to_slv(x : uint928_t) return std_logic_vector is
  variable rv : std_logic_vector(927 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint928_t(x : std_logic_vector) return uint928_t is
  variable rv : uint928_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int928_t_to_slv(x : int928_t) return std_logic_vector is
  variable rv : std_logic_vector(927 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int928_t(x : std_logic_vector) return int928_t is
  variable rv : int928_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint929_t_to_slv(x : uint929_t) return std_logic_vector is
  variable rv : std_logic_vector(928 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint929_t(x : std_logic_vector) return uint929_t is
  variable rv : uint929_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int929_t_to_slv(x : int929_t) return std_logic_vector is
  variable rv : std_logic_vector(928 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int929_t(x : std_logic_vector) return int929_t is
  variable rv : int929_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint930_t_to_slv(x : uint930_t) return std_logic_vector is
  variable rv : std_logic_vector(929 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint930_t(x : std_logic_vector) return uint930_t is
  variable rv : uint930_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int930_t_to_slv(x : int930_t) return std_logic_vector is
  variable rv : std_logic_vector(929 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int930_t(x : std_logic_vector) return int930_t is
  variable rv : int930_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint931_t_to_slv(x : uint931_t) return std_logic_vector is
  variable rv : std_logic_vector(930 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint931_t(x : std_logic_vector) return uint931_t is
  variable rv : uint931_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int931_t_to_slv(x : int931_t) return std_logic_vector is
  variable rv : std_logic_vector(930 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int931_t(x : std_logic_vector) return int931_t is
  variable rv : int931_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint932_t_to_slv(x : uint932_t) return std_logic_vector is
  variable rv : std_logic_vector(931 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint932_t(x : std_logic_vector) return uint932_t is
  variable rv : uint932_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int932_t_to_slv(x : int932_t) return std_logic_vector is
  variable rv : std_logic_vector(931 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int932_t(x : std_logic_vector) return int932_t is
  variable rv : int932_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint933_t_to_slv(x : uint933_t) return std_logic_vector is
  variable rv : std_logic_vector(932 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint933_t(x : std_logic_vector) return uint933_t is
  variable rv : uint933_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int933_t_to_slv(x : int933_t) return std_logic_vector is
  variable rv : std_logic_vector(932 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int933_t(x : std_logic_vector) return int933_t is
  variable rv : int933_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint934_t_to_slv(x : uint934_t) return std_logic_vector is
  variable rv : std_logic_vector(933 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint934_t(x : std_logic_vector) return uint934_t is
  variable rv : uint934_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int934_t_to_slv(x : int934_t) return std_logic_vector is
  variable rv : std_logic_vector(933 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int934_t(x : std_logic_vector) return int934_t is
  variable rv : int934_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint935_t_to_slv(x : uint935_t) return std_logic_vector is
  variable rv : std_logic_vector(934 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint935_t(x : std_logic_vector) return uint935_t is
  variable rv : uint935_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int935_t_to_slv(x : int935_t) return std_logic_vector is
  variable rv : std_logic_vector(934 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int935_t(x : std_logic_vector) return int935_t is
  variable rv : int935_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint936_t_to_slv(x : uint936_t) return std_logic_vector is
  variable rv : std_logic_vector(935 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint936_t(x : std_logic_vector) return uint936_t is
  variable rv : uint936_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int936_t_to_slv(x : int936_t) return std_logic_vector is
  variable rv : std_logic_vector(935 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int936_t(x : std_logic_vector) return int936_t is
  variable rv : int936_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint937_t_to_slv(x : uint937_t) return std_logic_vector is
  variable rv : std_logic_vector(936 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint937_t(x : std_logic_vector) return uint937_t is
  variable rv : uint937_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int937_t_to_slv(x : int937_t) return std_logic_vector is
  variable rv : std_logic_vector(936 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int937_t(x : std_logic_vector) return int937_t is
  variable rv : int937_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint938_t_to_slv(x : uint938_t) return std_logic_vector is
  variable rv : std_logic_vector(937 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint938_t(x : std_logic_vector) return uint938_t is
  variable rv : uint938_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int938_t_to_slv(x : int938_t) return std_logic_vector is
  variable rv : std_logic_vector(937 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int938_t(x : std_logic_vector) return int938_t is
  variable rv : int938_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint939_t_to_slv(x : uint939_t) return std_logic_vector is
  variable rv : std_logic_vector(938 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint939_t(x : std_logic_vector) return uint939_t is
  variable rv : uint939_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int939_t_to_slv(x : int939_t) return std_logic_vector is
  variable rv : std_logic_vector(938 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int939_t(x : std_logic_vector) return int939_t is
  variable rv : int939_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint940_t_to_slv(x : uint940_t) return std_logic_vector is
  variable rv : std_logic_vector(939 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint940_t(x : std_logic_vector) return uint940_t is
  variable rv : uint940_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int940_t_to_slv(x : int940_t) return std_logic_vector is
  variable rv : std_logic_vector(939 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int940_t(x : std_logic_vector) return int940_t is
  variable rv : int940_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint941_t_to_slv(x : uint941_t) return std_logic_vector is
  variable rv : std_logic_vector(940 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint941_t(x : std_logic_vector) return uint941_t is
  variable rv : uint941_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int941_t_to_slv(x : int941_t) return std_logic_vector is
  variable rv : std_logic_vector(940 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int941_t(x : std_logic_vector) return int941_t is
  variable rv : int941_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint942_t_to_slv(x : uint942_t) return std_logic_vector is
  variable rv : std_logic_vector(941 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint942_t(x : std_logic_vector) return uint942_t is
  variable rv : uint942_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int942_t_to_slv(x : int942_t) return std_logic_vector is
  variable rv : std_logic_vector(941 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int942_t(x : std_logic_vector) return int942_t is
  variable rv : int942_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint943_t_to_slv(x : uint943_t) return std_logic_vector is
  variable rv : std_logic_vector(942 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint943_t(x : std_logic_vector) return uint943_t is
  variable rv : uint943_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int943_t_to_slv(x : int943_t) return std_logic_vector is
  variable rv : std_logic_vector(942 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int943_t(x : std_logic_vector) return int943_t is
  variable rv : int943_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint944_t_to_slv(x : uint944_t) return std_logic_vector is
  variable rv : std_logic_vector(943 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint944_t(x : std_logic_vector) return uint944_t is
  variable rv : uint944_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int944_t_to_slv(x : int944_t) return std_logic_vector is
  variable rv : std_logic_vector(943 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int944_t(x : std_logic_vector) return int944_t is
  variable rv : int944_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint945_t_to_slv(x : uint945_t) return std_logic_vector is
  variable rv : std_logic_vector(944 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint945_t(x : std_logic_vector) return uint945_t is
  variable rv : uint945_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int945_t_to_slv(x : int945_t) return std_logic_vector is
  variable rv : std_logic_vector(944 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int945_t(x : std_logic_vector) return int945_t is
  variable rv : int945_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint946_t_to_slv(x : uint946_t) return std_logic_vector is
  variable rv : std_logic_vector(945 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint946_t(x : std_logic_vector) return uint946_t is
  variable rv : uint946_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int946_t_to_slv(x : int946_t) return std_logic_vector is
  variable rv : std_logic_vector(945 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int946_t(x : std_logic_vector) return int946_t is
  variable rv : int946_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint947_t_to_slv(x : uint947_t) return std_logic_vector is
  variable rv : std_logic_vector(946 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint947_t(x : std_logic_vector) return uint947_t is
  variable rv : uint947_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int947_t_to_slv(x : int947_t) return std_logic_vector is
  variable rv : std_logic_vector(946 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int947_t(x : std_logic_vector) return int947_t is
  variable rv : int947_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint948_t_to_slv(x : uint948_t) return std_logic_vector is
  variable rv : std_logic_vector(947 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint948_t(x : std_logic_vector) return uint948_t is
  variable rv : uint948_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int948_t_to_slv(x : int948_t) return std_logic_vector is
  variable rv : std_logic_vector(947 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int948_t(x : std_logic_vector) return int948_t is
  variable rv : int948_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint949_t_to_slv(x : uint949_t) return std_logic_vector is
  variable rv : std_logic_vector(948 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint949_t(x : std_logic_vector) return uint949_t is
  variable rv : uint949_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int949_t_to_slv(x : int949_t) return std_logic_vector is
  variable rv : std_logic_vector(948 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int949_t(x : std_logic_vector) return int949_t is
  variable rv : int949_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint950_t_to_slv(x : uint950_t) return std_logic_vector is
  variable rv : std_logic_vector(949 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint950_t(x : std_logic_vector) return uint950_t is
  variable rv : uint950_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int950_t_to_slv(x : int950_t) return std_logic_vector is
  variable rv : std_logic_vector(949 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int950_t(x : std_logic_vector) return int950_t is
  variable rv : int950_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint951_t_to_slv(x : uint951_t) return std_logic_vector is
  variable rv : std_logic_vector(950 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint951_t(x : std_logic_vector) return uint951_t is
  variable rv : uint951_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int951_t_to_slv(x : int951_t) return std_logic_vector is
  variable rv : std_logic_vector(950 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int951_t(x : std_logic_vector) return int951_t is
  variable rv : int951_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint952_t_to_slv(x : uint952_t) return std_logic_vector is
  variable rv : std_logic_vector(951 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint952_t(x : std_logic_vector) return uint952_t is
  variable rv : uint952_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int952_t_to_slv(x : int952_t) return std_logic_vector is
  variable rv : std_logic_vector(951 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int952_t(x : std_logic_vector) return int952_t is
  variable rv : int952_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint953_t_to_slv(x : uint953_t) return std_logic_vector is
  variable rv : std_logic_vector(952 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint953_t(x : std_logic_vector) return uint953_t is
  variable rv : uint953_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int953_t_to_slv(x : int953_t) return std_logic_vector is
  variable rv : std_logic_vector(952 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int953_t(x : std_logic_vector) return int953_t is
  variable rv : int953_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint954_t_to_slv(x : uint954_t) return std_logic_vector is
  variable rv : std_logic_vector(953 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint954_t(x : std_logic_vector) return uint954_t is
  variable rv : uint954_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int954_t_to_slv(x : int954_t) return std_logic_vector is
  variable rv : std_logic_vector(953 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int954_t(x : std_logic_vector) return int954_t is
  variable rv : int954_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint955_t_to_slv(x : uint955_t) return std_logic_vector is
  variable rv : std_logic_vector(954 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint955_t(x : std_logic_vector) return uint955_t is
  variable rv : uint955_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int955_t_to_slv(x : int955_t) return std_logic_vector is
  variable rv : std_logic_vector(954 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int955_t(x : std_logic_vector) return int955_t is
  variable rv : int955_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint956_t_to_slv(x : uint956_t) return std_logic_vector is
  variable rv : std_logic_vector(955 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint956_t(x : std_logic_vector) return uint956_t is
  variable rv : uint956_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int956_t_to_slv(x : int956_t) return std_logic_vector is
  variable rv : std_logic_vector(955 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int956_t(x : std_logic_vector) return int956_t is
  variable rv : int956_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint957_t_to_slv(x : uint957_t) return std_logic_vector is
  variable rv : std_logic_vector(956 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint957_t(x : std_logic_vector) return uint957_t is
  variable rv : uint957_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int957_t_to_slv(x : int957_t) return std_logic_vector is
  variable rv : std_logic_vector(956 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int957_t(x : std_logic_vector) return int957_t is
  variable rv : int957_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint958_t_to_slv(x : uint958_t) return std_logic_vector is
  variable rv : std_logic_vector(957 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint958_t(x : std_logic_vector) return uint958_t is
  variable rv : uint958_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int958_t_to_slv(x : int958_t) return std_logic_vector is
  variable rv : std_logic_vector(957 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int958_t(x : std_logic_vector) return int958_t is
  variable rv : int958_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint959_t_to_slv(x : uint959_t) return std_logic_vector is
  variable rv : std_logic_vector(958 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint959_t(x : std_logic_vector) return uint959_t is
  variable rv : uint959_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int959_t_to_slv(x : int959_t) return std_logic_vector is
  variable rv : std_logic_vector(958 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int959_t(x : std_logic_vector) return int959_t is
  variable rv : int959_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint960_t_to_slv(x : uint960_t) return std_logic_vector is
  variable rv : std_logic_vector(959 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint960_t(x : std_logic_vector) return uint960_t is
  variable rv : uint960_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int960_t_to_slv(x : int960_t) return std_logic_vector is
  variable rv : std_logic_vector(959 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int960_t(x : std_logic_vector) return int960_t is
  variable rv : int960_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint961_t_to_slv(x : uint961_t) return std_logic_vector is
  variable rv : std_logic_vector(960 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint961_t(x : std_logic_vector) return uint961_t is
  variable rv : uint961_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int961_t_to_slv(x : int961_t) return std_logic_vector is
  variable rv : std_logic_vector(960 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int961_t(x : std_logic_vector) return int961_t is
  variable rv : int961_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint962_t_to_slv(x : uint962_t) return std_logic_vector is
  variable rv : std_logic_vector(961 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint962_t(x : std_logic_vector) return uint962_t is
  variable rv : uint962_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int962_t_to_slv(x : int962_t) return std_logic_vector is
  variable rv : std_logic_vector(961 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int962_t(x : std_logic_vector) return int962_t is
  variable rv : int962_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint963_t_to_slv(x : uint963_t) return std_logic_vector is
  variable rv : std_logic_vector(962 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint963_t(x : std_logic_vector) return uint963_t is
  variable rv : uint963_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int963_t_to_slv(x : int963_t) return std_logic_vector is
  variable rv : std_logic_vector(962 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int963_t(x : std_logic_vector) return int963_t is
  variable rv : int963_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint964_t_to_slv(x : uint964_t) return std_logic_vector is
  variable rv : std_logic_vector(963 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint964_t(x : std_logic_vector) return uint964_t is
  variable rv : uint964_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int964_t_to_slv(x : int964_t) return std_logic_vector is
  variable rv : std_logic_vector(963 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int964_t(x : std_logic_vector) return int964_t is
  variable rv : int964_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint965_t_to_slv(x : uint965_t) return std_logic_vector is
  variable rv : std_logic_vector(964 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint965_t(x : std_logic_vector) return uint965_t is
  variable rv : uint965_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int965_t_to_slv(x : int965_t) return std_logic_vector is
  variable rv : std_logic_vector(964 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int965_t(x : std_logic_vector) return int965_t is
  variable rv : int965_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint966_t_to_slv(x : uint966_t) return std_logic_vector is
  variable rv : std_logic_vector(965 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint966_t(x : std_logic_vector) return uint966_t is
  variable rv : uint966_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int966_t_to_slv(x : int966_t) return std_logic_vector is
  variable rv : std_logic_vector(965 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int966_t(x : std_logic_vector) return int966_t is
  variable rv : int966_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint967_t_to_slv(x : uint967_t) return std_logic_vector is
  variable rv : std_logic_vector(966 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint967_t(x : std_logic_vector) return uint967_t is
  variable rv : uint967_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int967_t_to_slv(x : int967_t) return std_logic_vector is
  variable rv : std_logic_vector(966 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int967_t(x : std_logic_vector) return int967_t is
  variable rv : int967_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint968_t_to_slv(x : uint968_t) return std_logic_vector is
  variable rv : std_logic_vector(967 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint968_t(x : std_logic_vector) return uint968_t is
  variable rv : uint968_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int968_t_to_slv(x : int968_t) return std_logic_vector is
  variable rv : std_logic_vector(967 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int968_t(x : std_logic_vector) return int968_t is
  variable rv : int968_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint969_t_to_slv(x : uint969_t) return std_logic_vector is
  variable rv : std_logic_vector(968 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint969_t(x : std_logic_vector) return uint969_t is
  variable rv : uint969_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int969_t_to_slv(x : int969_t) return std_logic_vector is
  variable rv : std_logic_vector(968 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int969_t(x : std_logic_vector) return int969_t is
  variable rv : int969_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint970_t_to_slv(x : uint970_t) return std_logic_vector is
  variable rv : std_logic_vector(969 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint970_t(x : std_logic_vector) return uint970_t is
  variable rv : uint970_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int970_t_to_slv(x : int970_t) return std_logic_vector is
  variable rv : std_logic_vector(969 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int970_t(x : std_logic_vector) return int970_t is
  variable rv : int970_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint971_t_to_slv(x : uint971_t) return std_logic_vector is
  variable rv : std_logic_vector(970 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint971_t(x : std_logic_vector) return uint971_t is
  variable rv : uint971_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int971_t_to_slv(x : int971_t) return std_logic_vector is
  variable rv : std_logic_vector(970 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int971_t(x : std_logic_vector) return int971_t is
  variable rv : int971_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint972_t_to_slv(x : uint972_t) return std_logic_vector is
  variable rv : std_logic_vector(971 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint972_t(x : std_logic_vector) return uint972_t is
  variable rv : uint972_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int972_t_to_slv(x : int972_t) return std_logic_vector is
  variable rv : std_logic_vector(971 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int972_t(x : std_logic_vector) return int972_t is
  variable rv : int972_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint973_t_to_slv(x : uint973_t) return std_logic_vector is
  variable rv : std_logic_vector(972 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint973_t(x : std_logic_vector) return uint973_t is
  variable rv : uint973_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int973_t_to_slv(x : int973_t) return std_logic_vector is
  variable rv : std_logic_vector(972 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int973_t(x : std_logic_vector) return int973_t is
  variable rv : int973_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint974_t_to_slv(x : uint974_t) return std_logic_vector is
  variable rv : std_logic_vector(973 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint974_t(x : std_logic_vector) return uint974_t is
  variable rv : uint974_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int974_t_to_slv(x : int974_t) return std_logic_vector is
  variable rv : std_logic_vector(973 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int974_t(x : std_logic_vector) return int974_t is
  variable rv : int974_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint975_t_to_slv(x : uint975_t) return std_logic_vector is
  variable rv : std_logic_vector(974 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint975_t(x : std_logic_vector) return uint975_t is
  variable rv : uint975_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int975_t_to_slv(x : int975_t) return std_logic_vector is
  variable rv : std_logic_vector(974 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int975_t(x : std_logic_vector) return int975_t is
  variable rv : int975_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint976_t_to_slv(x : uint976_t) return std_logic_vector is
  variable rv : std_logic_vector(975 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint976_t(x : std_logic_vector) return uint976_t is
  variable rv : uint976_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int976_t_to_slv(x : int976_t) return std_logic_vector is
  variable rv : std_logic_vector(975 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int976_t(x : std_logic_vector) return int976_t is
  variable rv : int976_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint977_t_to_slv(x : uint977_t) return std_logic_vector is
  variable rv : std_logic_vector(976 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint977_t(x : std_logic_vector) return uint977_t is
  variable rv : uint977_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int977_t_to_slv(x : int977_t) return std_logic_vector is
  variable rv : std_logic_vector(976 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int977_t(x : std_logic_vector) return int977_t is
  variable rv : int977_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint978_t_to_slv(x : uint978_t) return std_logic_vector is
  variable rv : std_logic_vector(977 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint978_t(x : std_logic_vector) return uint978_t is
  variable rv : uint978_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int978_t_to_slv(x : int978_t) return std_logic_vector is
  variable rv : std_logic_vector(977 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int978_t(x : std_logic_vector) return int978_t is
  variable rv : int978_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint979_t_to_slv(x : uint979_t) return std_logic_vector is
  variable rv : std_logic_vector(978 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint979_t(x : std_logic_vector) return uint979_t is
  variable rv : uint979_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int979_t_to_slv(x : int979_t) return std_logic_vector is
  variable rv : std_logic_vector(978 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int979_t(x : std_logic_vector) return int979_t is
  variable rv : int979_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint980_t_to_slv(x : uint980_t) return std_logic_vector is
  variable rv : std_logic_vector(979 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint980_t(x : std_logic_vector) return uint980_t is
  variable rv : uint980_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int980_t_to_slv(x : int980_t) return std_logic_vector is
  variable rv : std_logic_vector(979 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int980_t(x : std_logic_vector) return int980_t is
  variable rv : int980_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint981_t_to_slv(x : uint981_t) return std_logic_vector is
  variable rv : std_logic_vector(980 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint981_t(x : std_logic_vector) return uint981_t is
  variable rv : uint981_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int981_t_to_slv(x : int981_t) return std_logic_vector is
  variable rv : std_logic_vector(980 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int981_t(x : std_logic_vector) return int981_t is
  variable rv : int981_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint982_t_to_slv(x : uint982_t) return std_logic_vector is
  variable rv : std_logic_vector(981 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint982_t(x : std_logic_vector) return uint982_t is
  variable rv : uint982_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int982_t_to_slv(x : int982_t) return std_logic_vector is
  variable rv : std_logic_vector(981 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int982_t(x : std_logic_vector) return int982_t is
  variable rv : int982_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint983_t_to_slv(x : uint983_t) return std_logic_vector is
  variable rv : std_logic_vector(982 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint983_t(x : std_logic_vector) return uint983_t is
  variable rv : uint983_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int983_t_to_slv(x : int983_t) return std_logic_vector is
  variable rv : std_logic_vector(982 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int983_t(x : std_logic_vector) return int983_t is
  variable rv : int983_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint984_t_to_slv(x : uint984_t) return std_logic_vector is
  variable rv : std_logic_vector(983 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint984_t(x : std_logic_vector) return uint984_t is
  variable rv : uint984_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int984_t_to_slv(x : int984_t) return std_logic_vector is
  variable rv : std_logic_vector(983 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int984_t(x : std_logic_vector) return int984_t is
  variable rv : int984_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint985_t_to_slv(x : uint985_t) return std_logic_vector is
  variable rv : std_logic_vector(984 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint985_t(x : std_logic_vector) return uint985_t is
  variable rv : uint985_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int985_t_to_slv(x : int985_t) return std_logic_vector is
  variable rv : std_logic_vector(984 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int985_t(x : std_logic_vector) return int985_t is
  variable rv : int985_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint986_t_to_slv(x : uint986_t) return std_logic_vector is
  variable rv : std_logic_vector(985 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint986_t(x : std_logic_vector) return uint986_t is
  variable rv : uint986_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int986_t_to_slv(x : int986_t) return std_logic_vector is
  variable rv : std_logic_vector(985 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int986_t(x : std_logic_vector) return int986_t is
  variable rv : int986_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint987_t_to_slv(x : uint987_t) return std_logic_vector is
  variable rv : std_logic_vector(986 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint987_t(x : std_logic_vector) return uint987_t is
  variable rv : uint987_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int987_t_to_slv(x : int987_t) return std_logic_vector is
  variable rv : std_logic_vector(986 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int987_t(x : std_logic_vector) return int987_t is
  variable rv : int987_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint988_t_to_slv(x : uint988_t) return std_logic_vector is
  variable rv : std_logic_vector(987 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint988_t(x : std_logic_vector) return uint988_t is
  variable rv : uint988_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int988_t_to_slv(x : int988_t) return std_logic_vector is
  variable rv : std_logic_vector(987 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int988_t(x : std_logic_vector) return int988_t is
  variable rv : int988_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint989_t_to_slv(x : uint989_t) return std_logic_vector is
  variable rv : std_logic_vector(988 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint989_t(x : std_logic_vector) return uint989_t is
  variable rv : uint989_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int989_t_to_slv(x : int989_t) return std_logic_vector is
  variable rv : std_logic_vector(988 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int989_t(x : std_logic_vector) return int989_t is
  variable rv : int989_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint990_t_to_slv(x : uint990_t) return std_logic_vector is
  variable rv : std_logic_vector(989 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint990_t(x : std_logic_vector) return uint990_t is
  variable rv : uint990_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int990_t_to_slv(x : int990_t) return std_logic_vector is
  variable rv : std_logic_vector(989 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int990_t(x : std_logic_vector) return int990_t is
  variable rv : int990_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint991_t_to_slv(x : uint991_t) return std_logic_vector is
  variable rv : std_logic_vector(990 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint991_t(x : std_logic_vector) return uint991_t is
  variable rv : uint991_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int991_t_to_slv(x : int991_t) return std_logic_vector is
  variable rv : std_logic_vector(990 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int991_t(x : std_logic_vector) return int991_t is
  variable rv : int991_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint992_t_to_slv(x : uint992_t) return std_logic_vector is
  variable rv : std_logic_vector(991 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint992_t(x : std_logic_vector) return uint992_t is
  variable rv : uint992_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int992_t_to_slv(x : int992_t) return std_logic_vector is
  variable rv : std_logic_vector(991 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int992_t(x : std_logic_vector) return int992_t is
  variable rv : int992_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint993_t_to_slv(x : uint993_t) return std_logic_vector is
  variable rv : std_logic_vector(992 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint993_t(x : std_logic_vector) return uint993_t is
  variable rv : uint993_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int993_t_to_slv(x : int993_t) return std_logic_vector is
  variable rv : std_logic_vector(992 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int993_t(x : std_logic_vector) return int993_t is
  variable rv : int993_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint994_t_to_slv(x : uint994_t) return std_logic_vector is
  variable rv : std_logic_vector(993 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint994_t(x : std_logic_vector) return uint994_t is
  variable rv : uint994_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int994_t_to_slv(x : int994_t) return std_logic_vector is
  variable rv : std_logic_vector(993 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int994_t(x : std_logic_vector) return int994_t is
  variable rv : int994_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint995_t_to_slv(x : uint995_t) return std_logic_vector is
  variable rv : std_logic_vector(994 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint995_t(x : std_logic_vector) return uint995_t is
  variable rv : uint995_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int995_t_to_slv(x : int995_t) return std_logic_vector is
  variable rv : std_logic_vector(994 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int995_t(x : std_logic_vector) return int995_t is
  variable rv : int995_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint996_t_to_slv(x : uint996_t) return std_logic_vector is
  variable rv : std_logic_vector(995 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint996_t(x : std_logic_vector) return uint996_t is
  variable rv : uint996_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int996_t_to_slv(x : int996_t) return std_logic_vector is
  variable rv : std_logic_vector(995 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int996_t(x : std_logic_vector) return int996_t is
  variable rv : int996_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint997_t_to_slv(x : uint997_t) return std_logic_vector is
  variable rv : std_logic_vector(996 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint997_t(x : std_logic_vector) return uint997_t is
  variable rv : uint997_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int997_t_to_slv(x : int997_t) return std_logic_vector is
  variable rv : std_logic_vector(996 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int997_t(x : std_logic_vector) return int997_t is
  variable rv : int997_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint998_t_to_slv(x : uint998_t) return std_logic_vector is
  variable rv : std_logic_vector(997 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint998_t(x : std_logic_vector) return uint998_t is
  variable rv : uint998_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int998_t_to_slv(x : int998_t) return std_logic_vector is
  variable rv : std_logic_vector(997 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int998_t(x : std_logic_vector) return int998_t is
  variable rv : int998_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint999_t_to_slv(x : uint999_t) return std_logic_vector is
  variable rv : std_logic_vector(998 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint999_t(x : std_logic_vector) return uint999_t is
  variable rv : uint999_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int999_t_to_slv(x : int999_t) return std_logic_vector is
  variable rv : std_logic_vector(998 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int999_t(x : std_logic_vector) return int999_t is
  variable rv : int999_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1000_t_to_slv(x : uint1000_t) return std_logic_vector is
  variable rv : std_logic_vector(999 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1000_t(x : std_logic_vector) return uint1000_t is
  variable rv : uint1000_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1000_t_to_slv(x : int1000_t) return std_logic_vector is
  variable rv : std_logic_vector(999 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1000_t(x : std_logic_vector) return int1000_t is
  variable rv : int1000_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1001_t_to_slv(x : uint1001_t) return std_logic_vector is
  variable rv : std_logic_vector(1000 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1001_t(x : std_logic_vector) return uint1001_t is
  variable rv : uint1001_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1001_t_to_slv(x : int1001_t) return std_logic_vector is
  variable rv : std_logic_vector(1000 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1001_t(x : std_logic_vector) return int1001_t is
  variable rv : int1001_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1002_t_to_slv(x : uint1002_t) return std_logic_vector is
  variable rv : std_logic_vector(1001 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1002_t(x : std_logic_vector) return uint1002_t is
  variable rv : uint1002_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1002_t_to_slv(x : int1002_t) return std_logic_vector is
  variable rv : std_logic_vector(1001 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1002_t(x : std_logic_vector) return int1002_t is
  variable rv : int1002_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1003_t_to_slv(x : uint1003_t) return std_logic_vector is
  variable rv : std_logic_vector(1002 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1003_t(x : std_logic_vector) return uint1003_t is
  variable rv : uint1003_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1003_t_to_slv(x : int1003_t) return std_logic_vector is
  variable rv : std_logic_vector(1002 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1003_t(x : std_logic_vector) return int1003_t is
  variable rv : int1003_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1004_t_to_slv(x : uint1004_t) return std_logic_vector is
  variable rv : std_logic_vector(1003 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1004_t(x : std_logic_vector) return uint1004_t is
  variable rv : uint1004_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1004_t_to_slv(x : int1004_t) return std_logic_vector is
  variable rv : std_logic_vector(1003 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1004_t(x : std_logic_vector) return int1004_t is
  variable rv : int1004_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1005_t_to_slv(x : uint1005_t) return std_logic_vector is
  variable rv : std_logic_vector(1004 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1005_t(x : std_logic_vector) return uint1005_t is
  variable rv : uint1005_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1005_t_to_slv(x : int1005_t) return std_logic_vector is
  variable rv : std_logic_vector(1004 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1005_t(x : std_logic_vector) return int1005_t is
  variable rv : int1005_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1006_t_to_slv(x : uint1006_t) return std_logic_vector is
  variable rv : std_logic_vector(1005 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1006_t(x : std_logic_vector) return uint1006_t is
  variable rv : uint1006_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1006_t_to_slv(x : int1006_t) return std_logic_vector is
  variable rv : std_logic_vector(1005 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1006_t(x : std_logic_vector) return int1006_t is
  variable rv : int1006_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1007_t_to_slv(x : uint1007_t) return std_logic_vector is
  variable rv : std_logic_vector(1006 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1007_t(x : std_logic_vector) return uint1007_t is
  variable rv : uint1007_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1007_t_to_slv(x : int1007_t) return std_logic_vector is
  variable rv : std_logic_vector(1006 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1007_t(x : std_logic_vector) return int1007_t is
  variable rv : int1007_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1008_t_to_slv(x : uint1008_t) return std_logic_vector is
  variable rv : std_logic_vector(1007 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1008_t(x : std_logic_vector) return uint1008_t is
  variable rv : uint1008_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1008_t_to_slv(x : int1008_t) return std_logic_vector is
  variable rv : std_logic_vector(1007 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1008_t(x : std_logic_vector) return int1008_t is
  variable rv : int1008_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1009_t_to_slv(x : uint1009_t) return std_logic_vector is
  variable rv : std_logic_vector(1008 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1009_t(x : std_logic_vector) return uint1009_t is
  variable rv : uint1009_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1009_t_to_slv(x : int1009_t) return std_logic_vector is
  variable rv : std_logic_vector(1008 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1009_t(x : std_logic_vector) return int1009_t is
  variable rv : int1009_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1010_t_to_slv(x : uint1010_t) return std_logic_vector is
  variable rv : std_logic_vector(1009 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1010_t(x : std_logic_vector) return uint1010_t is
  variable rv : uint1010_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1010_t_to_slv(x : int1010_t) return std_logic_vector is
  variable rv : std_logic_vector(1009 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1010_t(x : std_logic_vector) return int1010_t is
  variable rv : int1010_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1011_t_to_slv(x : uint1011_t) return std_logic_vector is
  variable rv : std_logic_vector(1010 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1011_t(x : std_logic_vector) return uint1011_t is
  variable rv : uint1011_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1011_t_to_slv(x : int1011_t) return std_logic_vector is
  variable rv : std_logic_vector(1010 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1011_t(x : std_logic_vector) return int1011_t is
  variable rv : int1011_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1012_t_to_slv(x : uint1012_t) return std_logic_vector is
  variable rv : std_logic_vector(1011 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1012_t(x : std_logic_vector) return uint1012_t is
  variable rv : uint1012_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1012_t_to_slv(x : int1012_t) return std_logic_vector is
  variable rv : std_logic_vector(1011 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1012_t(x : std_logic_vector) return int1012_t is
  variable rv : int1012_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1013_t_to_slv(x : uint1013_t) return std_logic_vector is
  variable rv : std_logic_vector(1012 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1013_t(x : std_logic_vector) return uint1013_t is
  variable rv : uint1013_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1013_t_to_slv(x : int1013_t) return std_logic_vector is
  variable rv : std_logic_vector(1012 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1013_t(x : std_logic_vector) return int1013_t is
  variable rv : int1013_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1014_t_to_slv(x : uint1014_t) return std_logic_vector is
  variable rv : std_logic_vector(1013 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1014_t(x : std_logic_vector) return uint1014_t is
  variable rv : uint1014_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1014_t_to_slv(x : int1014_t) return std_logic_vector is
  variable rv : std_logic_vector(1013 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1014_t(x : std_logic_vector) return int1014_t is
  variable rv : int1014_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1015_t_to_slv(x : uint1015_t) return std_logic_vector is
  variable rv : std_logic_vector(1014 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1015_t(x : std_logic_vector) return uint1015_t is
  variable rv : uint1015_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1015_t_to_slv(x : int1015_t) return std_logic_vector is
  variable rv : std_logic_vector(1014 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1015_t(x : std_logic_vector) return int1015_t is
  variable rv : int1015_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1016_t_to_slv(x : uint1016_t) return std_logic_vector is
  variable rv : std_logic_vector(1015 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1016_t(x : std_logic_vector) return uint1016_t is
  variable rv : uint1016_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1016_t_to_slv(x : int1016_t) return std_logic_vector is
  variable rv : std_logic_vector(1015 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1016_t(x : std_logic_vector) return int1016_t is
  variable rv : int1016_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1017_t_to_slv(x : uint1017_t) return std_logic_vector is
  variable rv : std_logic_vector(1016 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1017_t(x : std_logic_vector) return uint1017_t is
  variable rv : uint1017_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1017_t_to_slv(x : int1017_t) return std_logic_vector is
  variable rv : std_logic_vector(1016 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1017_t(x : std_logic_vector) return int1017_t is
  variable rv : int1017_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1018_t_to_slv(x : uint1018_t) return std_logic_vector is
  variable rv : std_logic_vector(1017 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1018_t(x : std_logic_vector) return uint1018_t is
  variable rv : uint1018_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1018_t_to_slv(x : int1018_t) return std_logic_vector is
  variable rv : std_logic_vector(1017 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1018_t(x : std_logic_vector) return int1018_t is
  variable rv : int1018_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1019_t_to_slv(x : uint1019_t) return std_logic_vector is
  variable rv : std_logic_vector(1018 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1019_t(x : std_logic_vector) return uint1019_t is
  variable rv : uint1019_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1019_t_to_slv(x : int1019_t) return std_logic_vector is
  variable rv : std_logic_vector(1018 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1019_t(x : std_logic_vector) return int1019_t is
  variable rv : int1019_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1020_t_to_slv(x : uint1020_t) return std_logic_vector is
  variable rv : std_logic_vector(1019 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1020_t(x : std_logic_vector) return uint1020_t is
  variable rv : uint1020_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1020_t_to_slv(x : int1020_t) return std_logic_vector is
  variable rv : std_logic_vector(1019 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1020_t(x : std_logic_vector) return int1020_t is
  variable rv : int1020_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1021_t_to_slv(x : uint1021_t) return std_logic_vector is
  variable rv : std_logic_vector(1020 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1021_t(x : std_logic_vector) return uint1021_t is
  variable rv : uint1021_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1021_t_to_slv(x : int1021_t) return std_logic_vector is
  variable rv : std_logic_vector(1020 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1021_t(x : std_logic_vector) return int1021_t is
  variable rv : int1021_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1022_t_to_slv(x : uint1022_t) return std_logic_vector is
  variable rv : std_logic_vector(1021 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1022_t(x : std_logic_vector) return uint1022_t is
  variable rv : uint1022_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1022_t_to_slv(x : int1022_t) return std_logic_vector is
  variable rv : std_logic_vector(1021 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1022_t(x : std_logic_vector) return int1022_t is
  variable rv : int1022_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1023_t_to_slv(x : uint1023_t) return std_logic_vector is
  variable rv : std_logic_vector(1022 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1023_t(x : std_logic_vector) return uint1023_t is
  variable rv : uint1023_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1023_t_to_slv(x : int1023_t) return std_logic_vector is
  variable rv : std_logic_vector(1022 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1023_t(x : std_logic_vector) return int1023_t is
  variable rv : int1023_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1024_t_to_slv(x : uint1024_t) return std_logic_vector is
  variable rv : std_logic_vector(1023 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1024_t(x : std_logic_vector) return uint1024_t is
  variable rv : uint1024_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1024_t_to_slv(x : int1024_t) return std_logic_vector is
  variable rv : std_logic_vector(1023 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1024_t(x : std_logic_vector) return int1024_t is
  variable rv : int1024_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1025_t_to_slv(x : uint1025_t) return std_logic_vector is
  variable rv : std_logic_vector(1024 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1025_t(x : std_logic_vector) return uint1025_t is
  variable rv : uint1025_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1025_t_to_slv(x : int1025_t) return std_logic_vector is
  variable rv : std_logic_vector(1024 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1025_t(x : std_logic_vector) return int1025_t is
  variable rv : int1025_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1026_t_to_slv(x : uint1026_t) return std_logic_vector is
  variable rv : std_logic_vector(1025 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1026_t(x : std_logic_vector) return uint1026_t is
  variable rv : uint1026_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1026_t_to_slv(x : int1026_t) return std_logic_vector is
  variable rv : std_logic_vector(1025 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1026_t(x : std_logic_vector) return int1026_t is
  variable rv : int1026_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1027_t_to_slv(x : uint1027_t) return std_logic_vector is
  variable rv : std_logic_vector(1026 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1027_t(x : std_logic_vector) return uint1027_t is
  variable rv : uint1027_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1027_t_to_slv(x : int1027_t) return std_logic_vector is
  variable rv : std_logic_vector(1026 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1027_t(x : std_logic_vector) return int1027_t is
  variable rv : int1027_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1028_t_to_slv(x : uint1028_t) return std_logic_vector is
  variable rv : std_logic_vector(1027 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1028_t(x : std_logic_vector) return uint1028_t is
  variable rv : uint1028_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1028_t_to_slv(x : int1028_t) return std_logic_vector is
  variable rv : std_logic_vector(1027 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1028_t(x : std_logic_vector) return int1028_t is
  variable rv : int1028_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1029_t_to_slv(x : uint1029_t) return std_logic_vector is
  variable rv : std_logic_vector(1028 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1029_t(x : std_logic_vector) return uint1029_t is
  variable rv : uint1029_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1029_t_to_slv(x : int1029_t) return std_logic_vector is
  variable rv : std_logic_vector(1028 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1029_t(x : std_logic_vector) return int1029_t is
  variable rv : int1029_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1030_t_to_slv(x : uint1030_t) return std_logic_vector is
  variable rv : std_logic_vector(1029 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1030_t(x : std_logic_vector) return uint1030_t is
  variable rv : uint1030_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1030_t_to_slv(x : int1030_t) return std_logic_vector is
  variable rv : std_logic_vector(1029 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1030_t(x : std_logic_vector) return int1030_t is
  variable rv : int1030_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1031_t_to_slv(x : uint1031_t) return std_logic_vector is
  variable rv : std_logic_vector(1030 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1031_t(x : std_logic_vector) return uint1031_t is
  variable rv : uint1031_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1031_t_to_slv(x : int1031_t) return std_logic_vector is
  variable rv : std_logic_vector(1030 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1031_t(x : std_logic_vector) return int1031_t is
  variable rv : int1031_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1032_t_to_slv(x : uint1032_t) return std_logic_vector is
  variable rv : std_logic_vector(1031 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1032_t(x : std_logic_vector) return uint1032_t is
  variable rv : uint1032_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1032_t_to_slv(x : int1032_t) return std_logic_vector is
  variable rv : std_logic_vector(1031 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1032_t(x : std_logic_vector) return int1032_t is
  variable rv : int1032_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1033_t_to_slv(x : uint1033_t) return std_logic_vector is
  variable rv : std_logic_vector(1032 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1033_t(x : std_logic_vector) return uint1033_t is
  variable rv : uint1033_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1033_t_to_slv(x : int1033_t) return std_logic_vector is
  variable rv : std_logic_vector(1032 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1033_t(x : std_logic_vector) return int1033_t is
  variable rv : int1033_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1034_t_to_slv(x : uint1034_t) return std_logic_vector is
  variable rv : std_logic_vector(1033 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1034_t(x : std_logic_vector) return uint1034_t is
  variable rv : uint1034_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1034_t_to_slv(x : int1034_t) return std_logic_vector is
  variable rv : std_logic_vector(1033 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1034_t(x : std_logic_vector) return int1034_t is
  variable rv : int1034_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1035_t_to_slv(x : uint1035_t) return std_logic_vector is
  variable rv : std_logic_vector(1034 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1035_t(x : std_logic_vector) return uint1035_t is
  variable rv : uint1035_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1035_t_to_slv(x : int1035_t) return std_logic_vector is
  variable rv : std_logic_vector(1034 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1035_t(x : std_logic_vector) return int1035_t is
  variable rv : int1035_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1036_t_to_slv(x : uint1036_t) return std_logic_vector is
  variable rv : std_logic_vector(1035 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1036_t(x : std_logic_vector) return uint1036_t is
  variable rv : uint1036_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1036_t_to_slv(x : int1036_t) return std_logic_vector is
  variable rv : std_logic_vector(1035 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1036_t(x : std_logic_vector) return int1036_t is
  variable rv : int1036_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1037_t_to_slv(x : uint1037_t) return std_logic_vector is
  variable rv : std_logic_vector(1036 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1037_t(x : std_logic_vector) return uint1037_t is
  variable rv : uint1037_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1037_t_to_slv(x : int1037_t) return std_logic_vector is
  variable rv : std_logic_vector(1036 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1037_t(x : std_logic_vector) return int1037_t is
  variable rv : int1037_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1038_t_to_slv(x : uint1038_t) return std_logic_vector is
  variable rv : std_logic_vector(1037 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1038_t(x : std_logic_vector) return uint1038_t is
  variable rv : uint1038_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1038_t_to_slv(x : int1038_t) return std_logic_vector is
  variable rv : std_logic_vector(1037 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1038_t(x : std_logic_vector) return int1038_t is
  variable rv : int1038_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1039_t_to_slv(x : uint1039_t) return std_logic_vector is
  variable rv : std_logic_vector(1038 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1039_t(x : std_logic_vector) return uint1039_t is
  variable rv : uint1039_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1039_t_to_slv(x : int1039_t) return std_logic_vector is
  variable rv : std_logic_vector(1038 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1039_t(x : std_logic_vector) return int1039_t is
  variable rv : int1039_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1040_t_to_slv(x : uint1040_t) return std_logic_vector is
  variable rv : std_logic_vector(1039 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1040_t(x : std_logic_vector) return uint1040_t is
  variable rv : uint1040_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1040_t_to_slv(x : int1040_t) return std_logic_vector is
  variable rv : std_logic_vector(1039 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1040_t(x : std_logic_vector) return int1040_t is
  variable rv : int1040_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1041_t_to_slv(x : uint1041_t) return std_logic_vector is
  variable rv : std_logic_vector(1040 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1041_t(x : std_logic_vector) return uint1041_t is
  variable rv : uint1041_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1041_t_to_slv(x : int1041_t) return std_logic_vector is
  variable rv : std_logic_vector(1040 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1041_t(x : std_logic_vector) return int1041_t is
  variable rv : int1041_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1042_t_to_slv(x : uint1042_t) return std_logic_vector is
  variable rv : std_logic_vector(1041 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1042_t(x : std_logic_vector) return uint1042_t is
  variable rv : uint1042_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1042_t_to_slv(x : int1042_t) return std_logic_vector is
  variable rv : std_logic_vector(1041 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1042_t(x : std_logic_vector) return int1042_t is
  variable rv : int1042_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1043_t_to_slv(x : uint1043_t) return std_logic_vector is
  variable rv : std_logic_vector(1042 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1043_t(x : std_logic_vector) return uint1043_t is
  variable rv : uint1043_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1043_t_to_slv(x : int1043_t) return std_logic_vector is
  variable rv : std_logic_vector(1042 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1043_t(x : std_logic_vector) return int1043_t is
  variable rv : int1043_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1044_t_to_slv(x : uint1044_t) return std_logic_vector is
  variable rv : std_logic_vector(1043 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1044_t(x : std_logic_vector) return uint1044_t is
  variable rv : uint1044_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1044_t_to_slv(x : int1044_t) return std_logic_vector is
  variable rv : std_logic_vector(1043 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1044_t(x : std_logic_vector) return int1044_t is
  variable rv : int1044_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1045_t_to_slv(x : uint1045_t) return std_logic_vector is
  variable rv : std_logic_vector(1044 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1045_t(x : std_logic_vector) return uint1045_t is
  variable rv : uint1045_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1045_t_to_slv(x : int1045_t) return std_logic_vector is
  variable rv : std_logic_vector(1044 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1045_t(x : std_logic_vector) return int1045_t is
  variable rv : int1045_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1046_t_to_slv(x : uint1046_t) return std_logic_vector is
  variable rv : std_logic_vector(1045 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1046_t(x : std_logic_vector) return uint1046_t is
  variable rv : uint1046_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1046_t_to_slv(x : int1046_t) return std_logic_vector is
  variable rv : std_logic_vector(1045 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1046_t(x : std_logic_vector) return int1046_t is
  variable rv : int1046_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1047_t_to_slv(x : uint1047_t) return std_logic_vector is
  variable rv : std_logic_vector(1046 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1047_t(x : std_logic_vector) return uint1047_t is
  variable rv : uint1047_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1047_t_to_slv(x : int1047_t) return std_logic_vector is
  variable rv : std_logic_vector(1046 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1047_t(x : std_logic_vector) return int1047_t is
  variable rv : int1047_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1048_t_to_slv(x : uint1048_t) return std_logic_vector is
  variable rv : std_logic_vector(1047 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1048_t(x : std_logic_vector) return uint1048_t is
  variable rv : uint1048_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1048_t_to_slv(x : int1048_t) return std_logic_vector is
  variable rv : std_logic_vector(1047 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1048_t(x : std_logic_vector) return int1048_t is
  variable rv : int1048_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1049_t_to_slv(x : uint1049_t) return std_logic_vector is
  variable rv : std_logic_vector(1048 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1049_t(x : std_logic_vector) return uint1049_t is
  variable rv : uint1049_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1049_t_to_slv(x : int1049_t) return std_logic_vector is
  variable rv : std_logic_vector(1048 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1049_t(x : std_logic_vector) return int1049_t is
  variable rv : int1049_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1050_t_to_slv(x : uint1050_t) return std_logic_vector is
  variable rv : std_logic_vector(1049 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1050_t(x : std_logic_vector) return uint1050_t is
  variable rv : uint1050_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1050_t_to_slv(x : int1050_t) return std_logic_vector is
  variable rv : std_logic_vector(1049 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1050_t(x : std_logic_vector) return int1050_t is
  variable rv : int1050_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1051_t_to_slv(x : uint1051_t) return std_logic_vector is
  variable rv : std_logic_vector(1050 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1051_t(x : std_logic_vector) return uint1051_t is
  variable rv : uint1051_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1051_t_to_slv(x : int1051_t) return std_logic_vector is
  variable rv : std_logic_vector(1050 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1051_t(x : std_logic_vector) return int1051_t is
  variable rv : int1051_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1052_t_to_slv(x : uint1052_t) return std_logic_vector is
  variable rv : std_logic_vector(1051 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1052_t(x : std_logic_vector) return uint1052_t is
  variable rv : uint1052_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1052_t_to_slv(x : int1052_t) return std_logic_vector is
  variable rv : std_logic_vector(1051 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1052_t(x : std_logic_vector) return int1052_t is
  variable rv : int1052_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1053_t_to_slv(x : uint1053_t) return std_logic_vector is
  variable rv : std_logic_vector(1052 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1053_t(x : std_logic_vector) return uint1053_t is
  variable rv : uint1053_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1053_t_to_slv(x : int1053_t) return std_logic_vector is
  variable rv : std_logic_vector(1052 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1053_t(x : std_logic_vector) return int1053_t is
  variable rv : int1053_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1054_t_to_slv(x : uint1054_t) return std_logic_vector is
  variable rv : std_logic_vector(1053 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1054_t(x : std_logic_vector) return uint1054_t is
  variable rv : uint1054_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1054_t_to_slv(x : int1054_t) return std_logic_vector is
  variable rv : std_logic_vector(1053 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1054_t(x : std_logic_vector) return int1054_t is
  variable rv : int1054_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1055_t_to_slv(x : uint1055_t) return std_logic_vector is
  variable rv : std_logic_vector(1054 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1055_t(x : std_logic_vector) return uint1055_t is
  variable rv : uint1055_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1055_t_to_slv(x : int1055_t) return std_logic_vector is
  variable rv : std_logic_vector(1054 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1055_t(x : std_logic_vector) return int1055_t is
  variable rv : int1055_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1056_t_to_slv(x : uint1056_t) return std_logic_vector is
  variable rv : std_logic_vector(1055 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1056_t(x : std_logic_vector) return uint1056_t is
  variable rv : uint1056_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1056_t_to_slv(x : int1056_t) return std_logic_vector is
  variable rv : std_logic_vector(1055 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1056_t(x : std_logic_vector) return int1056_t is
  variable rv : int1056_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1057_t_to_slv(x : uint1057_t) return std_logic_vector is
  variable rv : std_logic_vector(1056 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1057_t(x : std_logic_vector) return uint1057_t is
  variable rv : uint1057_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1057_t_to_slv(x : int1057_t) return std_logic_vector is
  variable rv : std_logic_vector(1056 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1057_t(x : std_logic_vector) return int1057_t is
  variable rv : int1057_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1058_t_to_slv(x : uint1058_t) return std_logic_vector is
  variable rv : std_logic_vector(1057 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1058_t(x : std_logic_vector) return uint1058_t is
  variable rv : uint1058_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1058_t_to_slv(x : int1058_t) return std_logic_vector is
  variable rv : std_logic_vector(1057 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1058_t(x : std_logic_vector) return int1058_t is
  variable rv : int1058_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1059_t_to_slv(x : uint1059_t) return std_logic_vector is
  variable rv : std_logic_vector(1058 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1059_t(x : std_logic_vector) return uint1059_t is
  variable rv : uint1059_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1059_t_to_slv(x : int1059_t) return std_logic_vector is
  variable rv : std_logic_vector(1058 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1059_t(x : std_logic_vector) return int1059_t is
  variable rv : int1059_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1060_t_to_slv(x : uint1060_t) return std_logic_vector is
  variable rv : std_logic_vector(1059 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1060_t(x : std_logic_vector) return uint1060_t is
  variable rv : uint1060_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1060_t_to_slv(x : int1060_t) return std_logic_vector is
  variable rv : std_logic_vector(1059 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1060_t(x : std_logic_vector) return int1060_t is
  variable rv : int1060_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1061_t_to_slv(x : uint1061_t) return std_logic_vector is
  variable rv : std_logic_vector(1060 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1061_t(x : std_logic_vector) return uint1061_t is
  variable rv : uint1061_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1061_t_to_slv(x : int1061_t) return std_logic_vector is
  variable rv : std_logic_vector(1060 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1061_t(x : std_logic_vector) return int1061_t is
  variable rv : int1061_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1062_t_to_slv(x : uint1062_t) return std_logic_vector is
  variable rv : std_logic_vector(1061 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1062_t(x : std_logic_vector) return uint1062_t is
  variable rv : uint1062_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1062_t_to_slv(x : int1062_t) return std_logic_vector is
  variable rv : std_logic_vector(1061 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1062_t(x : std_logic_vector) return int1062_t is
  variable rv : int1062_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1063_t_to_slv(x : uint1063_t) return std_logic_vector is
  variable rv : std_logic_vector(1062 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1063_t(x : std_logic_vector) return uint1063_t is
  variable rv : uint1063_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1063_t_to_slv(x : int1063_t) return std_logic_vector is
  variable rv : std_logic_vector(1062 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1063_t(x : std_logic_vector) return int1063_t is
  variable rv : int1063_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1064_t_to_slv(x : uint1064_t) return std_logic_vector is
  variable rv : std_logic_vector(1063 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1064_t(x : std_logic_vector) return uint1064_t is
  variable rv : uint1064_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1064_t_to_slv(x : int1064_t) return std_logic_vector is
  variable rv : std_logic_vector(1063 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1064_t(x : std_logic_vector) return int1064_t is
  variable rv : int1064_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1065_t_to_slv(x : uint1065_t) return std_logic_vector is
  variable rv : std_logic_vector(1064 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1065_t(x : std_logic_vector) return uint1065_t is
  variable rv : uint1065_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1065_t_to_slv(x : int1065_t) return std_logic_vector is
  variable rv : std_logic_vector(1064 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1065_t(x : std_logic_vector) return int1065_t is
  variable rv : int1065_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1066_t_to_slv(x : uint1066_t) return std_logic_vector is
  variable rv : std_logic_vector(1065 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1066_t(x : std_logic_vector) return uint1066_t is
  variable rv : uint1066_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1066_t_to_slv(x : int1066_t) return std_logic_vector is
  variable rv : std_logic_vector(1065 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1066_t(x : std_logic_vector) return int1066_t is
  variable rv : int1066_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1067_t_to_slv(x : uint1067_t) return std_logic_vector is
  variable rv : std_logic_vector(1066 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1067_t(x : std_logic_vector) return uint1067_t is
  variable rv : uint1067_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1067_t_to_slv(x : int1067_t) return std_logic_vector is
  variable rv : std_logic_vector(1066 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1067_t(x : std_logic_vector) return int1067_t is
  variable rv : int1067_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1068_t_to_slv(x : uint1068_t) return std_logic_vector is
  variable rv : std_logic_vector(1067 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1068_t(x : std_logic_vector) return uint1068_t is
  variable rv : uint1068_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1068_t_to_slv(x : int1068_t) return std_logic_vector is
  variable rv : std_logic_vector(1067 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1068_t(x : std_logic_vector) return int1068_t is
  variable rv : int1068_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1069_t_to_slv(x : uint1069_t) return std_logic_vector is
  variable rv : std_logic_vector(1068 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1069_t(x : std_logic_vector) return uint1069_t is
  variable rv : uint1069_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1069_t_to_slv(x : int1069_t) return std_logic_vector is
  variable rv : std_logic_vector(1068 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1069_t(x : std_logic_vector) return int1069_t is
  variable rv : int1069_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1070_t_to_slv(x : uint1070_t) return std_logic_vector is
  variable rv : std_logic_vector(1069 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1070_t(x : std_logic_vector) return uint1070_t is
  variable rv : uint1070_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1070_t_to_slv(x : int1070_t) return std_logic_vector is
  variable rv : std_logic_vector(1069 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1070_t(x : std_logic_vector) return int1070_t is
  variable rv : int1070_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1071_t_to_slv(x : uint1071_t) return std_logic_vector is
  variable rv : std_logic_vector(1070 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1071_t(x : std_logic_vector) return uint1071_t is
  variable rv : uint1071_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1071_t_to_slv(x : int1071_t) return std_logic_vector is
  variable rv : std_logic_vector(1070 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1071_t(x : std_logic_vector) return int1071_t is
  variable rv : int1071_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1072_t_to_slv(x : uint1072_t) return std_logic_vector is
  variable rv : std_logic_vector(1071 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1072_t(x : std_logic_vector) return uint1072_t is
  variable rv : uint1072_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1072_t_to_slv(x : int1072_t) return std_logic_vector is
  variable rv : std_logic_vector(1071 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1072_t(x : std_logic_vector) return int1072_t is
  variable rv : int1072_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1073_t_to_slv(x : uint1073_t) return std_logic_vector is
  variable rv : std_logic_vector(1072 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1073_t(x : std_logic_vector) return uint1073_t is
  variable rv : uint1073_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1073_t_to_slv(x : int1073_t) return std_logic_vector is
  variable rv : std_logic_vector(1072 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1073_t(x : std_logic_vector) return int1073_t is
  variable rv : int1073_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1074_t_to_slv(x : uint1074_t) return std_logic_vector is
  variable rv : std_logic_vector(1073 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1074_t(x : std_logic_vector) return uint1074_t is
  variable rv : uint1074_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1074_t_to_slv(x : int1074_t) return std_logic_vector is
  variable rv : std_logic_vector(1073 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1074_t(x : std_logic_vector) return int1074_t is
  variable rv : int1074_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1075_t_to_slv(x : uint1075_t) return std_logic_vector is
  variable rv : std_logic_vector(1074 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1075_t(x : std_logic_vector) return uint1075_t is
  variable rv : uint1075_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1075_t_to_slv(x : int1075_t) return std_logic_vector is
  variable rv : std_logic_vector(1074 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1075_t(x : std_logic_vector) return int1075_t is
  variable rv : int1075_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1076_t_to_slv(x : uint1076_t) return std_logic_vector is
  variable rv : std_logic_vector(1075 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1076_t(x : std_logic_vector) return uint1076_t is
  variable rv : uint1076_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1076_t_to_slv(x : int1076_t) return std_logic_vector is
  variable rv : std_logic_vector(1075 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1076_t(x : std_logic_vector) return int1076_t is
  variable rv : int1076_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1077_t_to_slv(x : uint1077_t) return std_logic_vector is
  variable rv : std_logic_vector(1076 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1077_t(x : std_logic_vector) return uint1077_t is
  variable rv : uint1077_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1077_t_to_slv(x : int1077_t) return std_logic_vector is
  variable rv : std_logic_vector(1076 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1077_t(x : std_logic_vector) return int1077_t is
  variable rv : int1077_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1078_t_to_slv(x : uint1078_t) return std_logic_vector is
  variable rv : std_logic_vector(1077 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1078_t(x : std_logic_vector) return uint1078_t is
  variable rv : uint1078_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1078_t_to_slv(x : int1078_t) return std_logic_vector is
  variable rv : std_logic_vector(1077 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1078_t(x : std_logic_vector) return int1078_t is
  variable rv : int1078_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1079_t_to_slv(x : uint1079_t) return std_logic_vector is
  variable rv : std_logic_vector(1078 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1079_t(x : std_logic_vector) return uint1079_t is
  variable rv : uint1079_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1079_t_to_slv(x : int1079_t) return std_logic_vector is
  variable rv : std_logic_vector(1078 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1079_t(x : std_logic_vector) return int1079_t is
  variable rv : int1079_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1080_t_to_slv(x : uint1080_t) return std_logic_vector is
  variable rv : std_logic_vector(1079 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1080_t(x : std_logic_vector) return uint1080_t is
  variable rv : uint1080_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1080_t_to_slv(x : int1080_t) return std_logic_vector is
  variable rv : std_logic_vector(1079 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1080_t(x : std_logic_vector) return int1080_t is
  variable rv : int1080_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1081_t_to_slv(x : uint1081_t) return std_logic_vector is
  variable rv : std_logic_vector(1080 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1081_t(x : std_logic_vector) return uint1081_t is
  variable rv : uint1081_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1081_t_to_slv(x : int1081_t) return std_logic_vector is
  variable rv : std_logic_vector(1080 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1081_t(x : std_logic_vector) return int1081_t is
  variable rv : int1081_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1082_t_to_slv(x : uint1082_t) return std_logic_vector is
  variable rv : std_logic_vector(1081 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1082_t(x : std_logic_vector) return uint1082_t is
  variable rv : uint1082_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1082_t_to_slv(x : int1082_t) return std_logic_vector is
  variable rv : std_logic_vector(1081 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1082_t(x : std_logic_vector) return int1082_t is
  variable rv : int1082_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1083_t_to_slv(x : uint1083_t) return std_logic_vector is
  variable rv : std_logic_vector(1082 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1083_t(x : std_logic_vector) return uint1083_t is
  variable rv : uint1083_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1083_t_to_slv(x : int1083_t) return std_logic_vector is
  variable rv : std_logic_vector(1082 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1083_t(x : std_logic_vector) return int1083_t is
  variable rv : int1083_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1084_t_to_slv(x : uint1084_t) return std_logic_vector is
  variable rv : std_logic_vector(1083 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1084_t(x : std_logic_vector) return uint1084_t is
  variable rv : uint1084_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1084_t_to_slv(x : int1084_t) return std_logic_vector is
  variable rv : std_logic_vector(1083 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1084_t(x : std_logic_vector) return int1084_t is
  variable rv : int1084_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1085_t_to_slv(x : uint1085_t) return std_logic_vector is
  variable rv : std_logic_vector(1084 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1085_t(x : std_logic_vector) return uint1085_t is
  variable rv : uint1085_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1085_t_to_slv(x : int1085_t) return std_logic_vector is
  variable rv : std_logic_vector(1084 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1085_t(x : std_logic_vector) return int1085_t is
  variable rv : int1085_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1086_t_to_slv(x : uint1086_t) return std_logic_vector is
  variable rv : std_logic_vector(1085 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1086_t(x : std_logic_vector) return uint1086_t is
  variable rv : uint1086_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1086_t_to_slv(x : int1086_t) return std_logic_vector is
  variable rv : std_logic_vector(1085 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1086_t(x : std_logic_vector) return int1086_t is
  variable rv : int1086_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1087_t_to_slv(x : uint1087_t) return std_logic_vector is
  variable rv : std_logic_vector(1086 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1087_t(x : std_logic_vector) return uint1087_t is
  variable rv : uint1087_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1087_t_to_slv(x : int1087_t) return std_logic_vector is
  variable rv : std_logic_vector(1086 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1087_t(x : std_logic_vector) return int1087_t is
  variable rv : int1087_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1088_t_to_slv(x : uint1088_t) return std_logic_vector is
  variable rv : std_logic_vector(1087 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1088_t(x : std_logic_vector) return uint1088_t is
  variable rv : uint1088_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1088_t_to_slv(x : int1088_t) return std_logic_vector is
  variable rv : std_logic_vector(1087 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1088_t(x : std_logic_vector) return int1088_t is
  variable rv : int1088_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1089_t_to_slv(x : uint1089_t) return std_logic_vector is
  variable rv : std_logic_vector(1088 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1089_t(x : std_logic_vector) return uint1089_t is
  variable rv : uint1089_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1089_t_to_slv(x : int1089_t) return std_logic_vector is
  variable rv : std_logic_vector(1088 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1089_t(x : std_logic_vector) return int1089_t is
  variable rv : int1089_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1090_t_to_slv(x : uint1090_t) return std_logic_vector is
  variable rv : std_logic_vector(1089 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1090_t(x : std_logic_vector) return uint1090_t is
  variable rv : uint1090_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1090_t_to_slv(x : int1090_t) return std_logic_vector is
  variable rv : std_logic_vector(1089 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1090_t(x : std_logic_vector) return int1090_t is
  variable rv : int1090_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1091_t_to_slv(x : uint1091_t) return std_logic_vector is
  variable rv : std_logic_vector(1090 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1091_t(x : std_logic_vector) return uint1091_t is
  variable rv : uint1091_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1091_t_to_slv(x : int1091_t) return std_logic_vector is
  variable rv : std_logic_vector(1090 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1091_t(x : std_logic_vector) return int1091_t is
  variable rv : int1091_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1092_t_to_slv(x : uint1092_t) return std_logic_vector is
  variable rv : std_logic_vector(1091 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1092_t(x : std_logic_vector) return uint1092_t is
  variable rv : uint1092_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1092_t_to_slv(x : int1092_t) return std_logic_vector is
  variable rv : std_logic_vector(1091 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1092_t(x : std_logic_vector) return int1092_t is
  variable rv : int1092_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1093_t_to_slv(x : uint1093_t) return std_logic_vector is
  variable rv : std_logic_vector(1092 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1093_t(x : std_logic_vector) return uint1093_t is
  variable rv : uint1093_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1093_t_to_slv(x : int1093_t) return std_logic_vector is
  variable rv : std_logic_vector(1092 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1093_t(x : std_logic_vector) return int1093_t is
  variable rv : int1093_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1094_t_to_slv(x : uint1094_t) return std_logic_vector is
  variable rv : std_logic_vector(1093 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1094_t(x : std_logic_vector) return uint1094_t is
  variable rv : uint1094_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1094_t_to_slv(x : int1094_t) return std_logic_vector is
  variable rv : std_logic_vector(1093 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1094_t(x : std_logic_vector) return int1094_t is
  variable rv : int1094_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1095_t_to_slv(x : uint1095_t) return std_logic_vector is
  variable rv : std_logic_vector(1094 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1095_t(x : std_logic_vector) return uint1095_t is
  variable rv : uint1095_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1095_t_to_slv(x : int1095_t) return std_logic_vector is
  variable rv : std_logic_vector(1094 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1095_t(x : std_logic_vector) return int1095_t is
  variable rv : int1095_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1096_t_to_slv(x : uint1096_t) return std_logic_vector is
  variable rv : std_logic_vector(1095 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1096_t(x : std_logic_vector) return uint1096_t is
  variable rv : uint1096_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1096_t_to_slv(x : int1096_t) return std_logic_vector is
  variable rv : std_logic_vector(1095 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1096_t(x : std_logic_vector) return int1096_t is
  variable rv : int1096_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1097_t_to_slv(x : uint1097_t) return std_logic_vector is
  variable rv : std_logic_vector(1096 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1097_t(x : std_logic_vector) return uint1097_t is
  variable rv : uint1097_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1097_t_to_slv(x : int1097_t) return std_logic_vector is
  variable rv : std_logic_vector(1096 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1097_t(x : std_logic_vector) return int1097_t is
  variable rv : int1097_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1098_t_to_slv(x : uint1098_t) return std_logic_vector is
  variable rv : std_logic_vector(1097 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1098_t(x : std_logic_vector) return uint1098_t is
  variable rv : uint1098_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1098_t_to_slv(x : int1098_t) return std_logic_vector is
  variable rv : std_logic_vector(1097 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1098_t(x : std_logic_vector) return int1098_t is
  variable rv : int1098_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1099_t_to_slv(x : uint1099_t) return std_logic_vector is
  variable rv : std_logic_vector(1098 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1099_t(x : std_logic_vector) return uint1099_t is
  variable rv : uint1099_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1099_t_to_slv(x : int1099_t) return std_logic_vector is
  variable rv : std_logic_vector(1098 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1099_t(x : std_logic_vector) return int1099_t is
  variable rv : int1099_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1100_t_to_slv(x : uint1100_t) return std_logic_vector is
  variable rv : std_logic_vector(1099 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1100_t(x : std_logic_vector) return uint1100_t is
  variable rv : uint1100_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1100_t_to_slv(x : int1100_t) return std_logic_vector is
  variable rv : std_logic_vector(1099 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1100_t(x : std_logic_vector) return int1100_t is
  variable rv : int1100_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1101_t_to_slv(x : uint1101_t) return std_logic_vector is
  variable rv : std_logic_vector(1100 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1101_t(x : std_logic_vector) return uint1101_t is
  variable rv : uint1101_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1101_t_to_slv(x : int1101_t) return std_logic_vector is
  variable rv : std_logic_vector(1100 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1101_t(x : std_logic_vector) return int1101_t is
  variable rv : int1101_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1102_t_to_slv(x : uint1102_t) return std_logic_vector is
  variable rv : std_logic_vector(1101 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1102_t(x : std_logic_vector) return uint1102_t is
  variable rv : uint1102_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1102_t_to_slv(x : int1102_t) return std_logic_vector is
  variable rv : std_logic_vector(1101 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1102_t(x : std_logic_vector) return int1102_t is
  variable rv : int1102_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1103_t_to_slv(x : uint1103_t) return std_logic_vector is
  variable rv : std_logic_vector(1102 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1103_t(x : std_logic_vector) return uint1103_t is
  variable rv : uint1103_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1103_t_to_slv(x : int1103_t) return std_logic_vector is
  variable rv : std_logic_vector(1102 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1103_t(x : std_logic_vector) return int1103_t is
  variable rv : int1103_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1104_t_to_slv(x : uint1104_t) return std_logic_vector is
  variable rv : std_logic_vector(1103 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1104_t(x : std_logic_vector) return uint1104_t is
  variable rv : uint1104_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1104_t_to_slv(x : int1104_t) return std_logic_vector is
  variable rv : std_logic_vector(1103 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1104_t(x : std_logic_vector) return int1104_t is
  variable rv : int1104_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1105_t_to_slv(x : uint1105_t) return std_logic_vector is
  variable rv : std_logic_vector(1104 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1105_t(x : std_logic_vector) return uint1105_t is
  variable rv : uint1105_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1105_t_to_slv(x : int1105_t) return std_logic_vector is
  variable rv : std_logic_vector(1104 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1105_t(x : std_logic_vector) return int1105_t is
  variable rv : int1105_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1106_t_to_slv(x : uint1106_t) return std_logic_vector is
  variable rv : std_logic_vector(1105 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1106_t(x : std_logic_vector) return uint1106_t is
  variable rv : uint1106_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1106_t_to_slv(x : int1106_t) return std_logic_vector is
  variable rv : std_logic_vector(1105 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1106_t(x : std_logic_vector) return int1106_t is
  variable rv : int1106_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1107_t_to_slv(x : uint1107_t) return std_logic_vector is
  variable rv : std_logic_vector(1106 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1107_t(x : std_logic_vector) return uint1107_t is
  variable rv : uint1107_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1107_t_to_slv(x : int1107_t) return std_logic_vector is
  variable rv : std_logic_vector(1106 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1107_t(x : std_logic_vector) return int1107_t is
  variable rv : int1107_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1108_t_to_slv(x : uint1108_t) return std_logic_vector is
  variable rv : std_logic_vector(1107 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1108_t(x : std_logic_vector) return uint1108_t is
  variable rv : uint1108_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1108_t_to_slv(x : int1108_t) return std_logic_vector is
  variable rv : std_logic_vector(1107 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1108_t(x : std_logic_vector) return int1108_t is
  variable rv : int1108_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1109_t_to_slv(x : uint1109_t) return std_logic_vector is
  variable rv : std_logic_vector(1108 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1109_t(x : std_logic_vector) return uint1109_t is
  variable rv : uint1109_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1109_t_to_slv(x : int1109_t) return std_logic_vector is
  variable rv : std_logic_vector(1108 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1109_t(x : std_logic_vector) return int1109_t is
  variable rv : int1109_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1110_t_to_slv(x : uint1110_t) return std_logic_vector is
  variable rv : std_logic_vector(1109 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1110_t(x : std_logic_vector) return uint1110_t is
  variable rv : uint1110_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1110_t_to_slv(x : int1110_t) return std_logic_vector is
  variable rv : std_logic_vector(1109 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1110_t(x : std_logic_vector) return int1110_t is
  variable rv : int1110_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1111_t_to_slv(x : uint1111_t) return std_logic_vector is
  variable rv : std_logic_vector(1110 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1111_t(x : std_logic_vector) return uint1111_t is
  variable rv : uint1111_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1111_t_to_slv(x : int1111_t) return std_logic_vector is
  variable rv : std_logic_vector(1110 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1111_t(x : std_logic_vector) return int1111_t is
  variable rv : int1111_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1112_t_to_slv(x : uint1112_t) return std_logic_vector is
  variable rv : std_logic_vector(1111 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1112_t(x : std_logic_vector) return uint1112_t is
  variable rv : uint1112_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1112_t_to_slv(x : int1112_t) return std_logic_vector is
  variable rv : std_logic_vector(1111 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1112_t(x : std_logic_vector) return int1112_t is
  variable rv : int1112_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1113_t_to_slv(x : uint1113_t) return std_logic_vector is
  variable rv : std_logic_vector(1112 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1113_t(x : std_logic_vector) return uint1113_t is
  variable rv : uint1113_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1113_t_to_slv(x : int1113_t) return std_logic_vector is
  variable rv : std_logic_vector(1112 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1113_t(x : std_logic_vector) return int1113_t is
  variable rv : int1113_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1114_t_to_slv(x : uint1114_t) return std_logic_vector is
  variable rv : std_logic_vector(1113 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1114_t(x : std_logic_vector) return uint1114_t is
  variable rv : uint1114_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1114_t_to_slv(x : int1114_t) return std_logic_vector is
  variable rv : std_logic_vector(1113 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1114_t(x : std_logic_vector) return int1114_t is
  variable rv : int1114_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1115_t_to_slv(x : uint1115_t) return std_logic_vector is
  variable rv : std_logic_vector(1114 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1115_t(x : std_logic_vector) return uint1115_t is
  variable rv : uint1115_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1115_t_to_slv(x : int1115_t) return std_logic_vector is
  variable rv : std_logic_vector(1114 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1115_t(x : std_logic_vector) return int1115_t is
  variable rv : int1115_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1116_t_to_slv(x : uint1116_t) return std_logic_vector is
  variable rv : std_logic_vector(1115 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1116_t(x : std_logic_vector) return uint1116_t is
  variable rv : uint1116_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1116_t_to_slv(x : int1116_t) return std_logic_vector is
  variable rv : std_logic_vector(1115 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1116_t(x : std_logic_vector) return int1116_t is
  variable rv : int1116_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1117_t_to_slv(x : uint1117_t) return std_logic_vector is
  variable rv : std_logic_vector(1116 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1117_t(x : std_logic_vector) return uint1117_t is
  variable rv : uint1117_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1117_t_to_slv(x : int1117_t) return std_logic_vector is
  variable rv : std_logic_vector(1116 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1117_t(x : std_logic_vector) return int1117_t is
  variable rv : int1117_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1118_t_to_slv(x : uint1118_t) return std_logic_vector is
  variable rv : std_logic_vector(1117 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1118_t(x : std_logic_vector) return uint1118_t is
  variable rv : uint1118_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1118_t_to_slv(x : int1118_t) return std_logic_vector is
  variable rv : std_logic_vector(1117 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1118_t(x : std_logic_vector) return int1118_t is
  variable rv : int1118_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1119_t_to_slv(x : uint1119_t) return std_logic_vector is
  variable rv : std_logic_vector(1118 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1119_t(x : std_logic_vector) return uint1119_t is
  variable rv : uint1119_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1119_t_to_slv(x : int1119_t) return std_logic_vector is
  variable rv : std_logic_vector(1118 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1119_t(x : std_logic_vector) return int1119_t is
  variable rv : int1119_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1120_t_to_slv(x : uint1120_t) return std_logic_vector is
  variable rv : std_logic_vector(1119 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1120_t(x : std_logic_vector) return uint1120_t is
  variable rv : uint1120_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1120_t_to_slv(x : int1120_t) return std_logic_vector is
  variable rv : std_logic_vector(1119 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1120_t(x : std_logic_vector) return int1120_t is
  variable rv : int1120_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1121_t_to_slv(x : uint1121_t) return std_logic_vector is
  variable rv : std_logic_vector(1120 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1121_t(x : std_logic_vector) return uint1121_t is
  variable rv : uint1121_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1121_t_to_slv(x : int1121_t) return std_logic_vector is
  variable rv : std_logic_vector(1120 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1121_t(x : std_logic_vector) return int1121_t is
  variable rv : int1121_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1122_t_to_slv(x : uint1122_t) return std_logic_vector is
  variable rv : std_logic_vector(1121 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1122_t(x : std_logic_vector) return uint1122_t is
  variable rv : uint1122_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1122_t_to_slv(x : int1122_t) return std_logic_vector is
  variable rv : std_logic_vector(1121 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1122_t(x : std_logic_vector) return int1122_t is
  variable rv : int1122_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1123_t_to_slv(x : uint1123_t) return std_logic_vector is
  variable rv : std_logic_vector(1122 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1123_t(x : std_logic_vector) return uint1123_t is
  variable rv : uint1123_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1123_t_to_slv(x : int1123_t) return std_logic_vector is
  variable rv : std_logic_vector(1122 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1123_t(x : std_logic_vector) return int1123_t is
  variable rv : int1123_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1124_t_to_slv(x : uint1124_t) return std_logic_vector is
  variable rv : std_logic_vector(1123 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1124_t(x : std_logic_vector) return uint1124_t is
  variable rv : uint1124_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1124_t_to_slv(x : int1124_t) return std_logic_vector is
  variable rv : std_logic_vector(1123 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1124_t(x : std_logic_vector) return int1124_t is
  variable rv : int1124_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1125_t_to_slv(x : uint1125_t) return std_logic_vector is
  variable rv : std_logic_vector(1124 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1125_t(x : std_logic_vector) return uint1125_t is
  variable rv : uint1125_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1125_t_to_slv(x : int1125_t) return std_logic_vector is
  variable rv : std_logic_vector(1124 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1125_t(x : std_logic_vector) return int1125_t is
  variable rv : int1125_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1126_t_to_slv(x : uint1126_t) return std_logic_vector is
  variable rv : std_logic_vector(1125 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1126_t(x : std_logic_vector) return uint1126_t is
  variable rv : uint1126_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1126_t_to_slv(x : int1126_t) return std_logic_vector is
  variable rv : std_logic_vector(1125 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1126_t(x : std_logic_vector) return int1126_t is
  variable rv : int1126_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1127_t_to_slv(x : uint1127_t) return std_logic_vector is
  variable rv : std_logic_vector(1126 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1127_t(x : std_logic_vector) return uint1127_t is
  variable rv : uint1127_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1127_t_to_slv(x : int1127_t) return std_logic_vector is
  variable rv : std_logic_vector(1126 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1127_t(x : std_logic_vector) return int1127_t is
  variable rv : int1127_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1128_t_to_slv(x : uint1128_t) return std_logic_vector is
  variable rv : std_logic_vector(1127 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1128_t(x : std_logic_vector) return uint1128_t is
  variable rv : uint1128_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1128_t_to_slv(x : int1128_t) return std_logic_vector is
  variable rv : std_logic_vector(1127 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1128_t(x : std_logic_vector) return int1128_t is
  variable rv : int1128_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1129_t_to_slv(x : uint1129_t) return std_logic_vector is
  variable rv : std_logic_vector(1128 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1129_t(x : std_logic_vector) return uint1129_t is
  variable rv : uint1129_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1129_t_to_slv(x : int1129_t) return std_logic_vector is
  variable rv : std_logic_vector(1128 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1129_t(x : std_logic_vector) return int1129_t is
  variable rv : int1129_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1130_t_to_slv(x : uint1130_t) return std_logic_vector is
  variable rv : std_logic_vector(1129 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1130_t(x : std_logic_vector) return uint1130_t is
  variable rv : uint1130_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1130_t_to_slv(x : int1130_t) return std_logic_vector is
  variable rv : std_logic_vector(1129 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1130_t(x : std_logic_vector) return int1130_t is
  variable rv : int1130_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1131_t_to_slv(x : uint1131_t) return std_logic_vector is
  variable rv : std_logic_vector(1130 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1131_t(x : std_logic_vector) return uint1131_t is
  variable rv : uint1131_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1131_t_to_slv(x : int1131_t) return std_logic_vector is
  variable rv : std_logic_vector(1130 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1131_t(x : std_logic_vector) return int1131_t is
  variable rv : int1131_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1132_t_to_slv(x : uint1132_t) return std_logic_vector is
  variable rv : std_logic_vector(1131 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1132_t(x : std_logic_vector) return uint1132_t is
  variable rv : uint1132_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1132_t_to_slv(x : int1132_t) return std_logic_vector is
  variable rv : std_logic_vector(1131 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1132_t(x : std_logic_vector) return int1132_t is
  variable rv : int1132_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1133_t_to_slv(x : uint1133_t) return std_logic_vector is
  variable rv : std_logic_vector(1132 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1133_t(x : std_logic_vector) return uint1133_t is
  variable rv : uint1133_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1133_t_to_slv(x : int1133_t) return std_logic_vector is
  variable rv : std_logic_vector(1132 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1133_t(x : std_logic_vector) return int1133_t is
  variable rv : int1133_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1134_t_to_slv(x : uint1134_t) return std_logic_vector is
  variable rv : std_logic_vector(1133 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1134_t(x : std_logic_vector) return uint1134_t is
  variable rv : uint1134_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1134_t_to_slv(x : int1134_t) return std_logic_vector is
  variable rv : std_logic_vector(1133 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1134_t(x : std_logic_vector) return int1134_t is
  variable rv : int1134_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1135_t_to_slv(x : uint1135_t) return std_logic_vector is
  variable rv : std_logic_vector(1134 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1135_t(x : std_logic_vector) return uint1135_t is
  variable rv : uint1135_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1135_t_to_slv(x : int1135_t) return std_logic_vector is
  variable rv : std_logic_vector(1134 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1135_t(x : std_logic_vector) return int1135_t is
  variable rv : int1135_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1136_t_to_slv(x : uint1136_t) return std_logic_vector is
  variable rv : std_logic_vector(1135 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1136_t(x : std_logic_vector) return uint1136_t is
  variable rv : uint1136_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1136_t_to_slv(x : int1136_t) return std_logic_vector is
  variable rv : std_logic_vector(1135 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1136_t(x : std_logic_vector) return int1136_t is
  variable rv : int1136_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1137_t_to_slv(x : uint1137_t) return std_logic_vector is
  variable rv : std_logic_vector(1136 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1137_t(x : std_logic_vector) return uint1137_t is
  variable rv : uint1137_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1137_t_to_slv(x : int1137_t) return std_logic_vector is
  variable rv : std_logic_vector(1136 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1137_t(x : std_logic_vector) return int1137_t is
  variable rv : int1137_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1138_t_to_slv(x : uint1138_t) return std_logic_vector is
  variable rv : std_logic_vector(1137 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1138_t(x : std_logic_vector) return uint1138_t is
  variable rv : uint1138_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1138_t_to_slv(x : int1138_t) return std_logic_vector is
  variable rv : std_logic_vector(1137 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1138_t(x : std_logic_vector) return int1138_t is
  variable rv : int1138_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1139_t_to_slv(x : uint1139_t) return std_logic_vector is
  variable rv : std_logic_vector(1138 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1139_t(x : std_logic_vector) return uint1139_t is
  variable rv : uint1139_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1139_t_to_slv(x : int1139_t) return std_logic_vector is
  variable rv : std_logic_vector(1138 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1139_t(x : std_logic_vector) return int1139_t is
  variable rv : int1139_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1140_t_to_slv(x : uint1140_t) return std_logic_vector is
  variable rv : std_logic_vector(1139 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1140_t(x : std_logic_vector) return uint1140_t is
  variable rv : uint1140_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1140_t_to_slv(x : int1140_t) return std_logic_vector is
  variable rv : std_logic_vector(1139 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1140_t(x : std_logic_vector) return int1140_t is
  variable rv : int1140_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1141_t_to_slv(x : uint1141_t) return std_logic_vector is
  variable rv : std_logic_vector(1140 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1141_t(x : std_logic_vector) return uint1141_t is
  variable rv : uint1141_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1141_t_to_slv(x : int1141_t) return std_logic_vector is
  variable rv : std_logic_vector(1140 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1141_t(x : std_logic_vector) return int1141_t is
  variable rv : int1141_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1142_t_to_slv(x : uint1142_t) return std_logic_vector is
  variable rv : std_logic_vector(1141 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1142_t(x : std_logic_vector) return uint1142_t is
  variable rv : uint1142_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1142_t_to_slv(x : int1142_t) return std_logic_vector is
  variable rv : std_logic_vector(1141 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1142_t(x : std_logic_vector) return int1142_t is
  variable rv : int1142_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1143_t_to_slv(x : uint1143_t) return std_logic_vector is
  variable rv : std_logic_vector(1142 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1143_t(x : std_logic_vector) return uint1143_t is
  variable rv : uint1143_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1143_t_to_slv(x : int1143_t) return std_logic_vector is
  variable rv : std_logic_vector(1142 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1143_t(x : std_logic_vector) return int1143_t is
  variable rv : int1143_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1144_t_to_slv(x : uint1144_t) return std_logic_vector is
  variable rv : std_logic_vector(1143 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1144_t(x : std_logic_vector) return uint1144_t is
  variable rv : uint1144_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1144_t_to_slv(x : int1144_t) return std_logic_vector is
  variable rv : std_logic_vector(1143 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1144_t(x : std_logic_vector) return int1144_t is
  variable rv : int1144_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1145_t_to_slv(x : uint1145_t) return std_logic_vector is
  variable rv : std_logic_vector(1144 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1145_t(x : std_logic_vector) return uint1145_t is
  variable rv : uint1145_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1145_t_to_slv(x : int1145_t) return std_logic_vector is
  variable rv : std_logic_vector(1144 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1145_t(x : std_logic_vector) return int1145_t is
  variable rv : int1145_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1146_t_to_slv(x : uint1146_t) return std_logic_vector is
  variable rv : std_logic_vector(1145 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1146_t(x : std_logic_vector) return uint1146_t is
  variable rv : uint1146_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1146_t_to_slv(x : int1146_t) return std_logic_vector is
  variable rv : std_logic_vector(1145 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1146_t(x : std_logic_vector) return int1146_t is
  variable rv : int1146_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1147_t_to_slv(x : uint1147_t) return std_logic_vector is
  variable rv : std_logic_vector(1146 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1147_t(x : std_logic_vector) return uint1147_t is
  variable rv : uint1147_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1147_t_to_slv(x : int1147_t) return std_logic_vector is
  variable rv : std_logic_vector(1146 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1147_t(x : std_logic_vector) return int1147_t is
  variable rv : int1147_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1148_t_to_slv(x : uint1148_t) return std_logic_vector is
  variable rv : std_logic_vector(1147 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1148_t(x : std_logic_vector) return uint1148_t is
  variable rv : uint1148_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1148_t_to_slv(x : int1148_t) return std_logic_vector is
  variable rv : std_logic_vector(1147 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1148_t(x : std_logic_vector) return int1148_t is
  variable rv : int1148_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1149_t_to_slv(x : uint1149_t) return std_logic_vector is
  variable rv : std_logic_vector(1148 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1149_t(x : std_logic_vector) return uint1149_t is
  variable rv : uint1149_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1149_t_to_slv(x : int1149_t) return std_logic_vector is
  variable rv : std_logic_vector(1148 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1149_t(x : std_logic_vector) return int1149_t is
  variable rv : int1149_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1150_t_to_slv(x : uint1150_t) return std_logic_vector is
  variable rv : std_logic_vector(1149 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1150_t(x : std_logic_vector) return uint1150_t is
  variable rv : uint1150_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1150_t_to_slv(x : int1150_t) return std_logic_vector is
  variable rv : std_logic_vector(1149 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1150_t(x : std_logic_vector) return int1150_t is
  variable rv : int1150_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1151_t_to_slv(x : uint1151_t) return std_logic_vector is
  variable rv : std_logic_vector(1150 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1151_t(x : std_logic_vector) return uint1151_t is
  variable rv : uint1151_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1151_t_to_slv(x : int1151_t) return std_logic_vector is
  variable rv : std_logic_vector(1150 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1151_t(x : std_logic_vector) return int1151_t is
  variable rv : int1151_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1152_t_to_slv(x : uint1152_t) return std_logic_vector is
  variable rv : std_logic_vector(1151 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1152_t(x : std_logic_vector) return uint1152_t is
  variable rv : uint1152_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1152_t_to_slv(x : int1152_t) return std_logic_vector is
  variable rv : std_logic_vector(1151 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1152_t(x : std_logic_vector) return int1152_t is
  variable rv : int1152_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1153_t_to_slv(x : uint1153_t) return std_logic_vector is
  variable rv : std_logic_vector(1152 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1153_t(x : std_logic_vector) return uint1153_t is
  variable rv : uint1153_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1153_t_to_slv(x : int1153_t) return std_logic_vector is
  variable rv : std_logic_vector(1152 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1153_t(x : std_logic_vector) return int1153_t is
  variable rv : int1153_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1154_t_to_slv(x : uint1154_t) return std_logic_vector is
  variable rv : std_logic_vector(1153 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1154_t(x : std_logic_vector) return uint1154_t is
  variable rv : uint1154_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1154_t_to_slv(x : int1154_t) return std_logic_vector is
  variable rv : std_logic_vector(1153 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1154_t(x : std_logic_vector) return int1154_t is
  variable rv : int1154_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1155_t_to_slv(x : uint1155_t) return std_logic_vector is
  variable rv : std_logic_vector(1154 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1155_t(x : std_logic_vector) return uint1155_t is
  variable rv : uint1155_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1155_t_to_slv(x : int1155_t) return std_logic_vector is
  variable rv : std_logic_vector(1154 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1155_t(x : std_logic_vector) return int1155_t is
  variable rv : int1155_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1156_t_to_slv(x : uint1156_t) return std_logic_vector is
  variable rv : std_logic_vector(1155 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1156_t(x : std_logic_vector) return uint1156_t is
  variable rv : uint1156_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1156_t_to_slv(x : int1156_t) return std_logic_vector is
  variable rv : std_logic_vector(1155 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1156_t(x : std_logic_vector) return int1156_t is
  variable rv : int1156_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1157_t_to_slv(x : uint1157_t) return std_logic_vector is
  variable rv : std_logic_vector(1156 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1157_t(x : std_logic_vector) return uint1157_t is
  variable rv : uint1157_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1157_t_to_slv(x : int1157_t) return std_logic_vector is
  variable rv : std_logic_vector(1156 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1157_t(x : std_logic_vector) return int1157_t is
  variable rv : int1157_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1158_t_to_slv(x : uint1158_t) return std_logic_vector is
  variable rv : std_logic_vector(1157 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1158_t(x : std_logic_vector) return uint1158_t is
  variable rv : uint1158_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1158_t_to_slv(x : int1158_t) return std_logic_vector is
  variable rv : std_logic_vector(1157 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1158_t(x : std_logic_vector) return int1158_t is
  variable rv : int1158_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1159_t_to_slv(x : uint1159_t) return std_logic_vector is
  variable rv : std_logic_vector(1158 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1159_t(x : std_logic_vector) return uint1159_t is
  variable rv : uint1159_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1159_t_to_slv(x : int1159_t) return std_logic_vector is
  variable rv : std_logic_vector(1158 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1159_t(x : std_logic_vector) return int1159_t is
  variable rv : int1159_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1160_t_to_slv(x : uint1160_t) return std_logic_vector is
  variable rv : std_logic_vector(1159 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1160_t(x : std_logic_vector) return uint1160_t is
  variable rv : uint1160_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1160_t_to_slv(x : int1160_t) return std_logic_vector is
  variable rv : std_logic_vector(1159 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1160_t(x : std_logic_vector) return int1160_t is
  variable rv : int1160_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1161_t_to_slv(x : uint1161_t) return std_logic_vector is
  variable rv : std_logic_vector(1160 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1161_t(x : std_logic_vector) return uint1161_t is
  variable rv : uint1161_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1161_t_to_slv(x : int1161_t) return std_logic_vector is
  variable rv : std_logic_vector(1160 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1161_t(x : std_logic_vector) return int1161_t is
  variable rv : int1161_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1162_t_to_slv(x : uint1162_t) return std_logic_vector is
  variable rv : std_logic_vector(1161 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1162_t(x : std_logic_vector) return uint1162_t is
  variable rv : uint1162_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1162_t_to_slv(x : int1162_t) return std_logic_vector is
  variable rv : std_logic_vector(1161 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1162_t(x : std_logic_vector) return int1162_t is
  variable rv : int1162_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1163_t_to_slv(x : uint1163_t) return std_logic_vector is
  variable rv : std_logic_vector(1162 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1163_t(x : std_logic_vector) return uint1163_t is
  variable rv : uint1163_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1163_t_to_slv(x : int1163_t) return std_logic_vector is
  variable rv : std_logic_vector(1162 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1163_t(x : std_logic_vector) return int1163_t is
  variable rv : int1163_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1164_t_to_slv(x : uint1164_t) return std_logic_vector is
  variable rv : std_logic_vector(1163 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1164_t(x : std_logic_vector) return uint1164_t is
  variable rv : uint1164_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1164_t_to_slv(x : int1164_t) return std_logic_vector is
  variable rv : std_logic_vector(1163 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1164_t(x : std_logic_vector) return int1164_t is
  variable rv : int1164_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1165_t_to_slv(x : uint1165_t) return std_logic_vector is
  variable rv : std_logic_vector(1164 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1165_t(x : std_logic_vector) return uint1165_t is
  variable rv : uint1165_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1165_t_to_slv(x : int1165_t) return std_logic_vector is
  variable rv : std_logic_vector(1164 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1165_t(x : std_logic_vector) return int1165_t is
  variable rv : int1165_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1166_t_to_slv(x : uint1166_t) return std_logic_vector is
  variable rv : std_logic_vector(1165 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1166_t(x : std_logic_vector) return uint1166_t is
  variable rv : uint1166_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1166_t_to_slv(x : int1166_t) return std_logic_vector is
  variable rv : std_logic_vector(1165 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1166_t(x : std_logic_vector) return int1166_t is
  variable rv : int1166_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1167_t_to_slv(x : uint1167_t) return std_logic_vector is
  variable rv : std_logic_vector(1166 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1167_t(x : std_logic_vector) return uint1167_t is
  variable rv : uint1167_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1167_t_to_slv(x : int1167_t) return std_logic_vector is
  variable rv : std_logic_vector(1166 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1167_t(x : std_logic_vector) return int1167_t is
  variable rv : int1167_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1168_t_to_slv(x : uint1168_t) return std_logic_vector is
  variable rv : std_logic_vector(1167 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1168_t(x : std_logic_vector) return uint1168_t is
  variable rv : uint1168_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1168_t_to_slv(x : int1168_t) return std_logic_vector is
  variable rv : std_logic_vector(1167 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1168_t(x : std_logic_vector) return int1168_t is
  variable rv : int1168_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1169_t_to_slv(x : uint1169_t) return std_logic_vector is
  variable rv : std_logic_vector(1168 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1169_t(x : std_logic_vector) return uint1169_t is
  variable rv : uint1169_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1169_t_to_slv(x : int1169_t) return std_logic_vector is
  variable rv : std_logic_vector(1168 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1169_t(x : std_logic_vector) return int1169_t is
  variable rv : int1169_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1170_t_to_slv(x : uint1170_t) return std_logic_vector is
  variable rv : std_logic_vector(1169 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1170_t(x : std_logic_vector) return uint1170_t is
  variable rv : uint1170_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1170_t_to_slv(x : int1170_t) return std_logic_vector is
  variable rv : std_logic_vector(1169 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1170_t(x : std_logic_vector) return int1170_t is
  variable rv : int1170_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1171_t_to_slv(x : uint1171_t) return std_logic_vector is
  variable rv : std_logic_vector(1170 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1171_t(x : std_logic_vector) return uint1171_t is
  variable rv : uint1171_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1171_t_to_slv(x : int1171_t) return std_logic_vector is
  variable rv : std_logic_vector(1170 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1171_t(x : std_logic_vector) return int1171_t is
  variable rv : int1171_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1172_t_to_slv(x : uint1172_t) return std_logic_vector is
  variable rv : std_logic_vector(1171 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1172_t(x : std_logic_vector) return uint1172_t is
  variable rv : uint1172_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1172_t_to_slv(x : int1172_t) return std_logic_vector is
  variable rv : std_logic_vector(1171 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1172_t(x : std_logic_vector) return int1172_t is
  variable rv : int1172_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1173_t_to_slv(x : uint1173_t) return std_logic_vector is
  variable rv : std_logic_vector(1172 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1173_t(x : std_logic_vector) return uint1173_t is
  variable rv : uint1173_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1173_t_to_slv(x : int1173_t) return std_logic_vector is
  variable rv : std_logic_vector(1172 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1173_t(x : std_logic_vector) return int1173_t is
  variable rv : int1173_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1174_t_to_slv(x : uint1174_t) return std_logic_vector is
  variable rv : std_logic_vector(1173 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1174_t(x : std_logic_vector) return uint1174_t is
  variable rv : uint1174_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1174_t_to_slv(x : int1174_t) return std_logic_vector is
  variable rv : std_logic_vector(1173 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1174_t(x : std_logic_vector) return int1174_t is
  variable rv : int1174_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1175_t_to_slv(x : uint1175_t) return std_logic_vector is
  variable rv : std_logic_vector(1174 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1175_t(x : std_logic_vector) return uint1175_t is
  variable rv : uint1175_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1175_t_to_slv(x : int1175_t) return std_logic_vector is
  variable rv : std_logic_vector(1174 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1175_t(x : std_logic_vector) return int1175_t is
  variable rv : int1175_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1176_t_to_slv(x : uint1176_t) return std_logic_vector is
  variable rv : std_logic_vector(1175 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1176_t(x : std_logic_vector) return uint1176_t is
  variable rv : uint1176_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1176_t_to_slv(x : int1176_t) return std_logic_vector is
  variable rv : std_logic_vector(1175 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1176_t(x : std_logic_vector) return int1176_t is
  variable rv : int1176_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1177_t_to_slv(x : uint1177_t) return std_logic_vector is
  variable rv : std_logic_vector(1176 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1177_t(x : std_logic_vector) return uint1177_t is
  variable rv : uint1177_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1177_t_to_slv(x : int1177_t) return std_logic_vector is
  variable rv : std_logic_vector(1176 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1177_t(x : std_logic_vector) return int1177_t is
  variable rv : int1177_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1178_t_to_slv(x : uint1178_t) return std_logic_vector is
  variable rv : std_logic_vector(1177 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1178_t(x : std_logic_vector) return uint1178_t is
  variable rv : uint1178_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1178_t_to_slv(x : int1178_t) return std_logic_vector is
  variable rv : std_logic_vector(1177 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1178_t(x : std_logic_vector) return int1178_t is
  variable rv : int1178_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1179_t_to_slv(x : uint1179_t) return std_logic_vector is
  variable rv : std_logic_vector(1178 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1179_t(x : std_logic_vector) return uint1179_t is
  variable rv : uint1179_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1179_t_to_slv(x : int1179_t) return std_logic_vector is
  variable rv : std_logic_vector(1178 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1179_t(x : std_logic_vector) return int1179_t is
  variable rv : int1179_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1180_t_to_slv(x : uint1180_t) return std_logic_vector is
  variable rv : std_logic_vector(1179 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1180_t(x : std_logic_vector) return uint1180_t is
  variable rv : uint1180_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1180_t_to_slv(x : int1180_t) return std_logic_vector is
  variable rv : std_logic_vector(1179 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1180_t(x : std_logic_vector) return int1180_t is
  variable rv : int1180_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1181_t_to_slv(x : uint1181_t) return std_logic_vector is
  variable rv : std_logic_vector(1180 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1181_t(x : std_logic_vector) return uint1181_t is
  variable rv : uint1181_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1181_t_to_slv(x : int1181_t) return std_logic_vector is
  variable rv : std_logic_vector(1180 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1181_t(x : std_logic_vector) return int1181_t is
  variable rv : int1181_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1182_t_to_slv(x : uint1182_t) return std_logic_vector is
  variable rv : std_logic_vector(1181 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1182_t(x : std_logic_vector) return uint1182_t is
  variable rv : uint1182_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1182_t_to_slv(x : int1182_t) return std_logic_vector is
  variable rv : std_logic_vector(1181 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1182_t(x : std_logic_vector) return int1182_t is
  variable rv : int1182_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1183_t_to_slv(x : uint1183_t) return std_logic_vector is
  variable rv : std_logic_vector(1182 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1183_t(x : std_logic_vector) return uint1183_t is
  variable rv : uint1183_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1183_t_to_slv(x : int1183_t) return std_logic_vector is
  variable rv : std_logic_vector(1182 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1183_t(x : std_logic_vector) return int1183_t is
  variable rv : int1183_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1184_t_to_slv(x : uint1184_t) return std_logic_vector is
  variable rv : std_logic_vector(1183 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1184_t(x : std_logic_vector) return uint1184_t is
  variable rv : uint1184_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1184_t_to_slv(x : int1184_t) return std_logic_vector is
  variable rv : std_logic_vector(1183 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1184_t(x : std_logic_vector) return int1184_t is
  variable rv : int1184_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1185_t_to_slv(x : uint1185_t) return std_logic_vector is
  variable rv : std_logic_vector(1184 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1185_t(x : std_logic_vector) return uint1185_t is
  variable rv : uint1185_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1185_t_to_slv(x : int1185_t) return std_logic_vector is
  variable rv : std_logic_vector(1184 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1185_t(x : std_logic_vector) return int1185_t is
  variable rv : int1185_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1186_t_to_slv(x : uint1186_t) return std_logic_vector is
  variable rv : std_logic_vector(1185 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1186_t(x : std_logic_vector) return uint1186_t is
  variable rv : uint1186_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1186_t_to_slv(x : int1186_t) return std_logic_vector is
  variable rv : std_logic_vector(1185 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1186_t(x : std_logic_vector) return int1186_t is
  variable rv : int1186_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1187_t_to_slv(x : uint1187_t) return std_logic_vector is
  variable rv : std_logic_vector(1186 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1187_t(x : std_logic_vector) return uint1187_t is
  variable rv : uint1187_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1187_t_to_slv(x : int1187_t) return std_logic_vector is
  variable rv : std_logic_vector(1186 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1187_t(x : std_logic_vector) return int1187_t is
  variable rv : int1187_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1188_t_to_slv(x : uint1188_t) return std_logic_vector is
  variable rv : std_logic_vector(1187 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1188_t(x : std_logic_vector) return uint1188_t is
  variable rv : uint1188_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1188_t_to_slv(x : int1188_t) return std_logic_vector is
  variable rv : std_logic_vector(1187 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1188_t(x : std_logic_vector) return int1188_t is
  variable rv : int1188_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1189_t_to_slv(x : uint1189_t) return std_logic_vector is
  variable rv : std_logic_vector(1188 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1189_t(x : std_logic_vector) return uint1189_t is
  variable rv : uint1189_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1189_t_to_slv(x : int1189_t) return std_logic_vector is
  variable rv : std_logic_vector(1188 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1189_t(x : std_logic_vector) return int1189_t is
  variable rv : int1189_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1190_t_to_slv(x : uint1190_t) return std_logic_vector is
  variable rv : std_logic_vector(1189 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1190_t(x : std_logic_vector) return uint1190_t is
  variable rv : uint1190_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1190_t_to_slv(x : int1190_t) return std_logic_vector is
  variable rv : std_logic_vector(1189 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1190_t(x : std_logic_vector) return int1190_t is
  variable rv : int1190_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1191_t_to_slv(x : uint1191_t) return std_logic_vector is
  variable rv : std_logic_vector(1190 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1191_t(x : std_logic_vector) return uint1191_t is
  variable rv : uint1191_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1191_t_to_slv(x : int1191_t) return std_logic_vector is
  variable rv : std_logic_vector(1190 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1191_t(x : std_logic_vector) return int1191_t is
  variable rv : int1191_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1192_t_to_slv(x : uint1192_t) return std_logic_vector is
  variable rv : std_logic_vector(1191 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1192_t(x : std_logic_vector) return uint1192_t is
  variable rv : uint1192_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1192_t_to_slv(x : int1192_t) return std_logic_vector is
  variable rv : std_logic_vector(1191 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1192_t(x : std_logic_vector) return int1192_t is
  variable rv : int1192_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1193_t_to_slv(x : uint1193_t) return std_logic_vector is
  variable rv : std_logic_vector(1192 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1193_t(x : std_logic_vector) return uint1193_t is
  variable rv : uint1193_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1193_t_to_slv(x : int1193_t) return std_logic_vector is
  variable rv : std_logic_vector(1192 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1193_t(x : std_logic_vector) return int1193_t is
  variable rv : int1193_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1194_t_to_slv(x : uint1194_t) return std_logic_vector is
  variable rv : std_logic_vector(1193 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1194_t(x : std_logic_vector) return uint1194_t is
  variable rv : uint1194_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1194_t_to_slv(x : int1194_t) return std_logic_vector is
  variable rv : std_logic_vector(1193 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1194_t(x : std_logic_vector) return int1194_t is
  variable rv : int1194_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1195_t_to_slv(x : uint1195_t) return std_logic_vector is
  variable rv : std_logic_vector(1194 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1195_t(x : std_logic_vector) return uint1195_t is
  variable rv : uint1195_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1195_t_to_slv(x : int1195_t) return std_logic_vector is
  variable rv : std_logic_vector(1194 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1195_t(x : std_logic_vector) return int1195_t is
  variable rv : int1195_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1196_t_to_slv(x : uint1196_t) return std_logic_vector is
  variable rv : std_logic_vector(1195 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1196_t(x : std_logic_vector) return uint1196_t is
  variable rv : uint1196_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1196_t_to_slv(x : int1196_t) return std_logic_vector is
  variable rv : std_logic_vector(1195 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1196_t(x : std_logic_vector) return int1196_t is
  variable rv : int1196_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1197_t_to_slv(x : uint1197_t) return std_logic_vector is
  variable rv : std_logic_vector(1196 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1197_t(x : std_logic_vector) return uint1197_t is
  variable rv : uint1197_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1197_t_to_slv(x : int1197_t) return std_logic_vector is
  variable rv : std_logic_vector(1196 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1197_t(x : std_logic_vector) return int1197_t is
  variable rv : int1197_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1198_t_to_slv(x : uint1198_t) return std_logic_vector is
  variable rv : std_logic_vector(1197 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1198_t(x : std_logic_vector) return uint1198_t is
  variable rv : uint1198_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1198_t_to_slv(x : int1198_t) return std_logic_vector is
  variable rv : std_logic_vector(1197 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1198_t(x : std_logic_vector) return int1198_t is
  variable rv : int1198_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1199_t_to_slv(x : uint1199_t) return std_logic_vector is
  variable rv : std_logic_vector(1198 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1199_t(x : std_logic_vector) return uint1199_t is
  variable rv : uint1199_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1199_t_to_slv(x : int1199_t) return std_logic_vector is
  variable rv : std_logic_vector(1198 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1199_t(x : std_logic_vector) return int1199_t is
  variable rv : int1199_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1200_t_to_slv(x : uint1200_t) return std_logic_vector is
  variable rv : std_logic_vector(1199 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1200_t(x : std_logic_vector) return uint1200_t is
  variable rv : uint1200_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1200_t_to_slv(x : int1200_t) return std_logic_vector is
  variable rv : std_logic_vector(1199 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1200_t(x : std_logic_vector) return int1200_t is
  variable rv : int1200_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1201_t_to_slv(x : uint1201_t) return std_logic_vector is
  variable rv : std_logic_vector(1200 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1201_t(x : std_logic_vector) return uint1201_t is
  variable rv : uint1201_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1201_t_to_slv(x : int1201_t) return std_logic_vector is
  variable rv : std_logic_vector(1200 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1201_t(x : std_logic_vector) return int1201_t is
  variable rv : int1201_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1202_t_to_slv(x : uint1202_t) return std_logic_vector is
  variable rv : std_logic_vector(1201 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1202_t(x : std_logic_vector) return uint1202_t is
  variable rv : uint1202_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1202_t_to_slv(x : int1202_t) return std_logic_vector is
  variable rv : std_logic_vector(1201 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1202_t(x : std_logic_vector) return int1202_t is
  variable rv : int1202_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1203_t_to_slv(x : uint1203_t) return std_logic_vector is
  variable rv : std_logic_vector(1202 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1203_t(x : std_logic_vector) return uint1203_t is
  variable rv : uint1203_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1203_t_to_slv(x : int1203_t) return std_logic_vector is
  variable rv : std_logic_vector(1202 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1203_t(x : std_logic_vector) return int1203_t is
  variable rv : int1203_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1204_t_to_slv(x : uint1204_t) return std_logic_vector is
  variable rv : std_logic_vector(1203 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1204_t(x : std_logic_vector) return uint1204_t is
  variable rv : uint1204_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1204_t_to_slv(x : int1204_t) return std_logic_vector is
  variable rv : std_logic_vector(1203 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1204_t(x : std_logic_vector) return int1204_t is
  variable rv : int1204_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1205_t_to_slv(x : uint1205_t) return std_logic_vector is
  variable rv : std_logic_vector(1204 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1205_t(x : std_logic_vector) return uint1205_t is
  variable rv : uint1205_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1205_t_to_slv(x : int1205_t) return std_logic_vector is
  variable rv : std_logic_vector(1204 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1205_t(x : std_logic_vector) return int1205_t is
  variable rv : int1205_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1206_t_to_slv(x : uint1206_t) return std_logic_vector is
  variable rv : std_logic_vector(1205 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1206_t(x : std_logic_vector) return uint1206_t is
  variable rv : uint1206_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1206_t_to_slv(x : int1206_t) return std_logic_vector is
  variable rv : std_logic_vector(1205 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1206_t(x : std_logic_vector) return int1206_t is
  variable rv : int1206_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1207_t_to_slv(x : uint1207_t) return std_logic_vector is
  variable rv : std_logic_vector(1206 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1207_t(x : std_logic_vector) return uint1207_t is
  variable rv : uint1207_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1207_t_to_slv(x : int1207_t) return std_logic_vector is
  variable rv : std_logic_vector(1206 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1207_t(x : std_logic_vector) return int1207_t is
  variable rv : int1207_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1208_t_to_slv(x : uint1208_t) return std_logic_vector is
  variable rv : std_logic_vector(1207 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1208_t(x : std_logic_vector) return uint1208_t is
  variable rv : uint1208_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1208_t_to_slv(x : int1208_t) return std_logic_vector is
  variable rv : std_logic_vector(1207 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1208_t(x : std_logic_vector) return int1208_t is
  variable rv : int1208_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1209_t_to_slv(x : uint1209_t) return std_logic_vector is
  variable rv : std_logic_vector(1208 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1209_t(x : std_logic_vector) return uint1209_t is
  variable rv : uint1209_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1209_t_to_slv(x : int1209_t) return std_logic_vector is
  variable rv : std_logic_vector(1208 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1209_t(x : std_logic_vector) return int1209_t is
  variable rv : int1209_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1210_t_to_slv(x : uint1210_t) return std_logic_vector is
  variable rv : std_logic_vector(1209 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1210_t(x : std_logic_vector) return uint1210_t is
  variable rv : uint1210_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1210_t_to_slv(x : int1210_t) return std_logic_vector is
  variable rv : std_logic_vector(1209 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1210_t(x : std_logic_vector) return int1210_t is
  variable rv : int1210_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1211_t_to_slv(x : uint1211_t) return std_logic_vector is
  variable rv : std_logic_vector(1210 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1211_t(x : std_logic_vector) return uint1211_t is
  variable rv : uint1211_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1211_t_to_slv(x : int1211_t) return std_logic_vector is
  variable rv : std_logic_vector(1210 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1211_t(x : std_logic_vector) return int1211_t is
  variable rv : int1211_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1212_t_to_slv(x : uint1212_t) return std_logic_vector is
  variable rv : std_logic_vector(1211 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1212_t(x : std_logic_vector) return uint1212_t is
  variable rv : uint1212_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1212_t_to_slv(x : int1212_t) return std_logic_vector is
  variable rv : std_logic_vector(1211 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1212_t(x : std_logic_vector) return int1212_t is
  variable rv : int1212_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1213_t_to_slv(x : uint1213_t) return std_logic_vector is
  variable rv : std_logic_vector(1212 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1213_t(x : std_logic_vector) return uint1213_t is
  variable rv : uint1213_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1213_t_to_slv(x : int1213_t) return std_logic_vector is
  variable rv : std_logic_vector(1212 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1213_t(x : std_logic_vector) return int1213_t is
  variable rv : int1213_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1214_t_to_slv(x : uint1214_t) return std_logic_vector is
  variable rv : std_logic_vector(1213 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1214_t(x : std_logic_vector) return uint1214_t is
  variable rv : uint1214_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1214_t_to_slv(x : int1214_t) return std_logic_vector is
  variable rv : std_logic_vector(1213 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1214_t(x : std_logic_vector) return int1214_t is
  variable rv : int1214_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1215_t_to_slv(x : uint1215_t) return std_logic_vector is
  variable rv : std_logic_vector(1214 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1215_t(x : std_logic_vector) return uint1215_t is
  variable rv : uint1215_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1215_t_to_slv(x : int1215_t) return std_logic_vector is
  variable rv : std_logic_vector(1214 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1215_t(x : std_logic_vector) return int1215_t is
  variable rv : int1215_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1216_t_to_slv(x : uint1216_t) return std_logic_vector is
  variable rv : std_logic_vector(1215 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1216_t(x : std_logic_vector) return uint1216_t is
  variable rv : uint1216_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1216_t_to_slv(x : int1216_t) return std_logic_vector is
  variable rv : std_logic_vector(1215 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1216_t(x : std_logic_vector) return int1216_t is
  variable rv : int1216_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1217_t_to_slv(x : uint1217_t) return std_logic_vector is
  variable rv : std_logic_vector(1216 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1217_t(x : std_logic_vector) return uint1217_t is
  variable rv : uint1217_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1217_t_to_slv(x : int1217_t) return std_logic_vector is
  variable rv : std_logic_vector(1216 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1217_t(x : std_logic_vector) return int1217_t is
  variable rv : int1217_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1218_t_to_slv(x : uint1218_t) return std_logic_vector is
  variable rv : std_logic_vector(1217 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1218_t(x : std_logic_vector) return uint1218_t is
  variable rv : uint1218_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1218_t_to_slv(x : int1218_t) return std_logic_vector is
  variable rv : std_logic_vector(1217 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1218_t(x : std_logic_vector) return int1218_t is
  variable rv : int1218_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1219_t_to_slv(x : uint1219_t) return std_logic_vector is
  variable rv : std_logic_vector(1218 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1219_t(x : std_logic_vector) return uint1219_t is
  variable rv : uint1219_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1219_t_to_slv(x : int1219_t) return std_logic_vector is
  variable rv : std_logic_vector(1218 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1219_t(x : std_logic_vector) return int1219_t is
  variable rv : int1219_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1220_t_to_slv(x : uint1220_t) return std_logic_vector is
  variable rv : std_logic_vector(1219 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1220_t(x : std_logic_vector) return uint1220_t is
  variable rv : uint1220_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1220_t_to_slv(x : int1220_t) return std_logic_vector is
  variable rv : std_logic_vector(1219 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1220_t(x : std_logic_vector) return int1220_t is
  variable rv : int1220_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1221_t_to_slv(x : uint1221_t) return std_logic_vector is
  variable rv : std_logic_vector(1220 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1221_t(x : std_logic_vector) return uint1221_t is
  variable rv : uint1221_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1221_t_to_slv(x : int1221_t) return std_logic_vector is
  variable rv : std_logic_vector(1220 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1221_t(x : std_logic_vector) return int1221_t is
  variable rv : int1221_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1222_t_to_slv(x : uint1222_t) return std_logic_vector is
  variable rv : std_logic_vector(1221 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1222_t(x : std_logic_vector) return uint1222_t is
  variable rv : uint1222_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1222_t_to_slv(x : int1222_t) return std_logic_vector is
  variable rv : std_logic_vector(1221 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1222_t(x : std_logic_vector) return int1222_t is
  variable rv : int1222_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1223_t_to_slv(x : uint1223_t) return std_logic_vector is
  variable rv : std_logic_vector(1222 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1223_t(x : std_logic_vector) return uint1223_t is
  variable rv : uint1223_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1223_t_to_slv(x : int1223_t) return std_logic_vector is
  variable rv : std_logic_vector(1222 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1223_t(x : std_logic_vector) return int1223_t is
  variable rv : int1223_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1224_t_to_slv(x : uint1224_t) return std_logic_vector is
  variable rv : std_logic_vector(1223 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1224_t(x : std_logic_vector) return uint1224_t is
  variable rv : uint1224_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1224_t_to_slv(x : int1224_t) return std_logic_vector is
  variable rv : std_logic_vector(1223 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1224_t(x : std_logic_vector) return int1224_t is
  variable rv : int1224_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1225_t_to_slv(x : uint1225_t) return std_logic_vector is
  variable rv : std_logic_vector(1224 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1225_t(x : std_logic_vector) return uint1225_t is
  variable rv : uint1225_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1225_t_to_slv(x : int1225_t) return std_logic_vector is
  variable rv : std_logic_vector(1224 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1225_t(x : std_logic_vector) return int1225_t is
  variable rv : int1225_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1226_t_to_slv(x : uint1226_t) return std_logic_vector is
  variable rv : std_logic_vector(1225 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1226_t(x : std_logic_vector) return uint1226_t is
  variable rv : uint1226_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1226_t_to_slv(x : int1226_t) return std_logic_vector is
  variable rv : std_logic_vector(1225 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1226_t(x : std_logic_vector) return int1226_t is
  variable rv : int1226_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1227_t_to_slv(x : uint1227_t) return std_logic_vector is
  variable rv : std_logic_vector(1226 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1227_t(x : std_logic_vector) return uint1227_t is
  variable rv : uint1227_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1227_t_to_slv(x : int1227_t) return std_logic_vector is
  variable rv : std_logic_vector(1226 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1227_t(x : std_logic_vector) return int1227_t is
  variable rv : int1227_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1228_t_to_slv(x : uint1228_t) return std_logic_vector is
  variable rv : std_logic_vector(1227 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1228_t(x : std_logic_vector) return uint1228_t is
  variable rv : uint1228_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1228_t_to_slv(x : int1228_t) return std_logic_vector is
  variable rv : std_logic_vector(1227 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1228_t(x : std_logic_vector) return int1228_t is
  variable rv : int1228_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1229_t_to_slv(x : uint1229_t) return std_logic_vector is
  variable rv : std_logic_vector(1228 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1229_t(x : std_logic_vector) return uint1229_t is
  variable rv : uint1229_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1229_t_to_slv(x : int1229_t) return std_logic_vector is
  variable rv : std_logic_vector(1228 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1229_t(x : std_logic_vector) return int1229_t is
  variable rv : int1229_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1230_t_to_slv(x : uint1230_t) return std_logic_vector is
  variable rv : std_logic_vector(1229 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1230_t(x : std_logic_vector) return uint1230_t is
  variable rv : uint1230_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1230_t_to_slv(x : int1230_t) return std_logic_vector is
  variable rv : std_logic_vector(1229 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1230_t(x : std_logic_vector) return int1230_t is
  variable rv : int1230_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1231_t_to_slv(x : uint1231_t) return std_logic_vector is
  variable rv : std_logic_vector(1230 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1231_t(x : std_logic_vector) return uint1231_t is
  variable rv : uint1231_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1231_t_to_slv(x : int1231_t) return std_logic_vector is
  variable rv : std_logic_vector(1230 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1231_t(x : std_logic_vector) return int1231_t is
  variable rv : int1231_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1232_t_to_slv(x : uint1232_t) return std_logic_vector is
  variable rv : std_logic_vector(1231 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1232_t(x : std_logic_vector) return uint1232_t is
  variable rv : uint1232_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1232_t_to_slv(x : int1232_t) return std_logic_vector is
  variable rv : std_logic_vector(1231 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1232_t(x : std_logic_vector) return int1232_t is
  variable rv : int1232_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1233_t_to_slv(x : uint1233_t) return std_logic_vector is
  variable rv : std_logic_vector(1232 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1233_t(x : std_logic_vector) return uint1233_t is
  variable rv : uint1233_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1233_t_to_slv(x : int1233_t) return std_logic_vector is
  variable rv : std_logic_vector(1232 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1233_t(x : std_logic_vector) return int1233_t is
  variable rv : int1233_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1234_t_to_slv(x : uint1234_t) return std_logic_vector is
  variable rv : std_logic_vector(1233 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1234_t(x : std_logic_vector) return uint1234_t is
  variable rv : uint1234_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1234_t_to_slv(x : int1234_t) return std_logic_vector is
  variable rv : std_logic_vector(1233 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1234_t(x : std_logic_vector) return int1234_t is
  variable rv : int1234_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1235_t_to_slv(x : uint1235_t) return std_logic_vector is
  variable rv : std_logic_vector(1234 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1235_t(x : std_logic_vector) return uint1235_t is
  variable rv : uint1235_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1235_t_to_slv(x : int1235_t) return std_logic_vector is
  variable rv : std_logic_vector(1234 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1235_t(x : std_logic_vector) return int1235_t is
  variable rv : int1235_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1236_t_to_slv(x : uint1236_t) return std_logic_vector is
  variable rv : std_logic_vector(1235 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1236_t(x : std_logic_vector) return uint1236_t is
  variable rv : uint1236_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1236_t_to_slv(x : int1236_t) return std_logic_vector is
  variable rv : std_logic_vector(1235 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1236_t(x : std_logic_vector) return int1236_t is
  variable rv : int1236_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1237_t_to_slv(x : uint1237_t) return std_logic_vector is
  variable rv : std_logic_vector(1236 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1237_t(x : std_logic_vector) return uint1237_t is
  variable rv : uint1237_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1237_t_to_slv(x : int1237_t) return std_logic_vector is
  variable rv : std_logic_vector(1236 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1237_t(x : std_logic_vector) return int1237_t is
  variable rv : int1237_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1238_t_to_slv(x : uint1238_t) return std_logic_vector is
  variable rv : std_logic_vector(1237 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1238_t(x : std_logic_vector) return uint1238_t is
  variable rv : uint1238_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1238_t_to_slv(x : int1238_t) return std_logic_vector is
  variable rv : std_logic_vector(1237 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1238_t(x : std_logic_vector) return int1238_t is
  variable rv : int1238_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1239_t_to_slv(x : uint1239_t) return std_logic_vector is
  variable rv : std_logic_vector(1238 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1239_t(x : std_logic_vector) return uint1239_t is
  variable rv : uint1239_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1239_t_to_slv(x : int1239_t) return std_logic_vector is
  variable rv : std_logic_vector(1238 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1239_t(x : std_logic_vector) return int1239_t is
  variable rv : int1239_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1240_t_to_slv(x : uint1240_t) return std_logic_vector is
  variable rv : std_logic_vector(1239 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1240_t(x : std_logic_vector) return uint1240_t is
  variable rv : uint1240_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1240_t_to_slv(x : int1240_t) return std_logic_vector is
  variable rv : std_logic_vector(1239 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1240_t(x : std_logic_vector) return int1240_t is
  variable rv : int1240_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1241_t_to_slv(x : uint1241_t) return std_logic_vector is
  variable rv : std_logic_vector(1240 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1241_t(x : std_logic_vector) return uint1241_t is
  variable rv : uint1241_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1241_t_to_slv(x : int1241_t) return std_logic_vector is
  variable rv : std_logic_vector(1240 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1241_t(x : std_logic_vector) return int1241_t is
  variable rv : int1241_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1242_t_to_slv(x : uint1242_t) return std_logic_vector is
  variable rv : std_logic_vector(1241 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1242_t(x : std_logic_vector) return uint1242_t is
  variable rv : uint1242_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1242_t_to_slv(x : int1242_t) return std_logic_vector is
  variable rv : std_logic_vector(1241 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1242_t(x : std_logic_vector) return int1242_t is
  variable rv : int1242_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1243_t_to_slv(x : uint1243_t) return std_logic_vector is
  variable rv : std_logic_vector(1242 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1243_t(x : std_logic_vector) return uint1243_t is
  variable rv : uint1243_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1243_t_to_slv(x : int1243_t) return std_logic_vector is
  variable rv : std_logic_vector(1242 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1243_t(x : std_logic_vector) return int1243_t is
  variable rv : int1243_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1244_t_to_slv(x : uint1244_t) return std_logic_vector is
  variable rv : std_logic_vector(1243 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1244_t(x : std_logic_vector) return uint1244_t is
  variable rv : uint1244_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1244_t_to_slv(x : int1244_t) return std_logic_vector is
  variable rv : std_logic_vector(1243 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1244_t(x : std_logic_vector) return int1244_t is
  variable rv : int1244_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1245_t_to_slv(x : uint1245_t) return std_logic_vector is
  variable rv : std_logic_vector(1244 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1245_t(x : std_logic_vector) return uint1245_t is
  variable rv : uint1245_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1245_t_to_slv(x : int1245_t) return std_logic_vector is
  variable rv : std_logic_vector(1244 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1245_t(x : std_logic_vector) return int1245_t is
  variable rv : int1245_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1246_t_to_slv(x : uint1246_t) return std_logic_vector is
  variable rv : std_logic_vector(1245 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1246_t(x : std_logic_vector) return uint1246_t is
  variable rv : uint1246_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1246_t_to_slv(x : int1246_t) return std_logic_vector is
  variable rv : std_logic_vector(1245 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1246_t(x : std_logic_vector) return int1246_t is
  variable rv : int1246_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1247_t_to_slv(x : uint1247_t) return std_logic_vector is
  variable rv : std_logic_vector(1246 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1247_t(x : std_logic_vector) return uint1247_t is
  variable rv : uint1247_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1247_t_to_slv(x : int1247_t) return std_logic_vector is
  variable rv : std_logic_vector(1246 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1247_t(x : std_logic_vector) return int1247_t is
  variable rv : int1247_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1248_t_to_slv(x : uint1248_t) return std_logic_vector is
  variable rv : std_logic_vector(1247 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1248_t(x : std_logic_vector) return uint1248_t is
  variable rv : uint1248_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1248_t_to_slv(x : int1248_t) return std_logic_vector is
  variable rv : std_logic_vector(1247 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1248_t(x : std_logic_vector) return int1248_t is
  variable rv : int1248_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1249_t_to_slv(x : uint1249_t) return std_logic_vector is
  variable rv : std_logic_vector(1248 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1249_t(x : std_logic_vector) return uint1249_t is
  variable rv : uint1249_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1249_t_to_slv(x : int1249_t) return std_logic_vector is
  variable rv : std_logic_vector(1248 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1249_t(x : std_logic_vector) return int1249_t is
  variable rv : int1249_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1250_t_to_slv(x : uint1250_t) return std_logic_vector is
  variable rv : std_logic_vector(1249 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1250_t(x : std_logic_vector) return uint1250_t is
  variable rv : uint1250_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1250_t_to_slv(x : int1250_t) return std_logic_vector is
  variable rv : std_logic_vector(1249 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1250_t(x : std_logic_vector) return int1250_t is
  variable rv : int1250_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1251_t_to_slv(x : uint1251_t) return std_logic_vector is
  variable rv : std_logic_vector(1250 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1251_t(x : std_logic_vector) return uint1251_t is
  variable rv : uint1251_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1251_t_to_slv(x : int1251_t) return std_logic_vector is
  variable rv : std_logic_vector(1250 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1251_t(x : std_logic_vector) return int1251_t is
  variable rv : int1251_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1252_t_to_slv(x : uint1252_t) return std_logic_vector is
  variable rv : std_logic_vector(1251 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1252_t(x : std_logic_vector) return uint1252_t is
  variable rv : uint1252_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1252_t_to_slv(x : int1252_t) return std_logic_vector is
  variable rv : std_logic_vector(1251 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1252_t(x : std_logic_vector) return int1252_t is
  variable rv : int1252_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1253_t_to_slv(x : uint1253_t) return std_logic_vector is
  variable rv : std_logic_vector(1252 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1253_t(x : std_logic_vector) return uint1253_t is
  variable rv : uint1253_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1253_t_to_slv(x : int1253_t) return std_logic_vector is
  variable rv : std_logic_vector(1252 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1253_t(x : std_logic_vector) return int1253_t is
  variable rv : int1253_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1254_t_to_slv(x : uint1254_t) return std_logic_vector is
  variable rv : std_logic_vector(1253 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1254_t(x : std_logic_vector) return uint1254_t is
  variable rv : uint1254_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1254_t_to_slv(x : int1254_t) return std_logic_vector is
  variable rv : std_logic_vector(1253 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1254_t(x : std_logic_vector) return int1254_t is
  variable rv : int1254_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1255_t_to_slv(x : uint1255_t) return std_logic_vector is
  variable rv : std_logic_vector(1254 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1255_t(x : std_logic_vector) return uint1255_t is
  variable rv : uint1255_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1255_t_to_slv(x : int1255_t) return std_logic_vector is
  variable rv : std_logic_vector(1254 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1255_t(x : std_logic_vector) return int1255_t is
  variable rv : int1255_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1256_t_to_slv(x : uint1256_t) return std_logic_vector is
  variable rv : std_logic_vector(1255 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1256_t(x : std_logic_vector) return uint1256_t is
  variable rv : uint1256_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1256_t_to_slv(x : int1256_t) return std_logic_vector is
  variable rv : std_logic_vector(1255 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1256_t(x : std_logic_vector) return int1256_t is
  variable rv : int1256_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1257_t_to_slv(x : uint1257_t) return std_logic_vector is
  variable rv : std_logic_vector(1256 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1257_t(x : std_logic_vector) return uint1257_t is
  variable rv : uint1257_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1257_t_to_slv(x : int1257_t) return std_logic_vector is
  variable rv : std_logic_vector(1256 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1257_t(x : std_logic_vector) return int1257_t is
  variable rv : int1257_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1258_t_to_slv(x : uint1258_t) return std_logic_vector is
  variable rv : std_logic_vector(1257 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1258_t(x : std_logic_vector) return uint1258_t is
  variable rv : uint1258_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1258_t_to_slv(x : int1258_t) return std_logic_vector is
  variable rv : std_logic_vector(1257 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1258_t(x : std_logic_vector) return int1258_t is
  variable rv : int1258_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1259_t_to_slv(x : uint1259_t) return std_logic_vector is
  variable rv : std_logic_vector(1258 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1259_t(x : std_logic_vector) return uint1259_t is
  variable rv : uint1259_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1259_t_to_slv(x : int1259_t) return std_logic_vector is
  variable rv : std_logic_vector(1258 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1259_t(x : std_logic_vector) return int1259_t is
  variable rv : int1259_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1260_t_to_slv(x : uint1260_t) return std_logic_vector is
  variable rv : std_logic_vector(1259 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1260_t(x : std_logic_vector) return uint1260_t is
  variable rv : uint1260_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1260_t_to_slv(x : int1260_t) return std_logic_vector is
  variable rv : std_logic_vector(1259 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1260_t(x : std_logic_vector) return int1260_t is
  variable rv : int1260_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1261_t_to_slv(x : uint1261_t) return std_logic_vector is
  variable rv : std_logic_vector(1260 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1261_t(x : std_logic_vector) return uint1261_t is
  variable rv : uint1261_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1261_t_to_slv(x : int1261_t) return std_logic_vector is
  variable rv : std_logic_vector(1260 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1261_t(x : std_logic_vector) return int1261_t is
  variable rv : int1261_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1262_t_to_slv(x : uint1262_t) return std_logic_vector is
  variable rv : std_logic_vector(1261 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1262_t(x : std_logic_vector) return uint1262_t is
  variable rv : uint1262_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1262_t_to_slv(x : int1262_t) return std_logic_vector is
  variable rv : std_logic_vector(1261 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1262_t(x : std_logic_vector) return int1262_t is
  variable rv : int1262_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1263_t_to_slv(x : uint1263_t) return std_logic_vector is
  variable rv : std_logic_vector(1262 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1263_t(x : std_logic_vector) return uint1263_t is
  variable rv : uint1263_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1263_t_to_slv(x : int1263_t) return std_logic_vector is
  variable rv : std_logic_vector(1262 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1263_t(x : std_logic_vector) return int1263_t is
  variable rv : int1263_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1264_t_to_slv(x : uint1264_t) return std_logic_vector is
  variable rv : std_logic_vector(1263 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1264_t(x : std_logic_vector) return uint1264_t is
  variable rv : uint1264_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1264_t_to_slv(x : int1264_t) return std_logic_vector is
  variable rv : std_logic_vector(1263 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1264_t(x : std_logic_vector) return int1264_t is
  variable rv : int1264_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1265_t_to_slv(x : uint1265_t) return std_logic_vector is
  variable rv : std_logic_vector(1264 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1265_t(x : std_logic_vector) return uint1265_t is
  variable rv : uint1265_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1265_t_to_slv(x : int1265_t) return std_logic_vector is
  variable rv : std_logic_vector(1264 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1265_t(x : std_logic_vector) return int1265_t is
  variable rv : int1265_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1266_t_to_slv(x : uint1266_t) return std_logic_vector is
  variable rv : std_logic_vector(1265 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1266_t(x : std_logic_vector) return uint1266_t is
  variable rv : uint1266_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1266_t_to_slv(x : int1266_t) return std_logic_vector is
  variable rv : std_logic_vector(1265 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1266_t(x : std_logic_vector) return int1266_t is
  variable rv : int1266_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1267_t_to_slv(x : uint1267_t) return std_logic_vector is
  variable rv : std_logic_vector(1266 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1267_t(x : std_logic_vector) return uint1267_t is
  variable rv : uint1267_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1267_t_to_slv(x : int1267_t) return std_logic_vector is
  variable rv : std_logic_vector(1266 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1267_t(x : std_logic_vector) return int1267_t is
  variable rv : int1267_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1268_t_to_slv(x : uint1268_t) return std_logic_vector is
  variable rv : std_logic_vector(1267 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1268_t(x : std_logic_vector) return uint1268_t is
  variable rv : uint1268_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1268_t_to_slv(x : int1268_t) return std_logic_vector is
  variable rv : std_logic_vector(1267 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1268_t(x : std_logic_vector) return int1268_t is
  variable rv : int1268_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1269_t_to_slv(x : uint1269_t) return std_logic_vector is
  variable rv : std_logic_vector(1268 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1269_t(x : std_logic_vector) return uint1269_t is
  variable rv : uint1269_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1269_t_to_slv(x : int1269_t) return std_logic_vector is
  variable rv : std_logic_vector(1268 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1269_t(x : std_logic_vector) return int1269_t is
  variable rv : int1269_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1270_t_to_slv(x : uint1270_t) return std_logic_vector is
  variable rv : std_logic_vector(1269 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1270_t(x : std_logic_vector) return uint1270_t is
  variable rv : uint1270_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1270_t_to_slv(x : int1270_t) return std_logic_vector is
  variable rv : std_logic_vector(1269 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1270_t(x : std_logic_vector) return int1270_t is
  variable rv : int1270_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1271_t_to_slv(x : uint1271_t) return std_logic_vector is
  variable rv : std_logic_vector(1270 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1271_t(x : std_logic_vector) return uint1271_t is
  variable rv : uint1271_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1271_t_to_slv(x : int1271_t) return std_logic_vector is
  variable rv : std_logic_vector(1270 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1271_t(x : std_logic_vector) return int1271_t is
  variable rv : int1271_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1272_t_to_slv(x : uint1272_t) return std_logic_vector is
  variable rv : std_logic_vector(1271 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1272_t(x : std_logic_vector) return uint1272_t is
  variable rv : uint1272_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1272_t_to_slv(x : int1272_t) return std_logic_vector is
  variable rv : std_logic_vector(1271 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1272_t(x : std_logic_vector) return int1272_t is
  variable rv : int1272_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1273_t_to_slv(x : uint1273_t) return std_logic_vector is
  variable rv : std_logic_vector(1272 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1273_t(x : std_logic_vector) return uint1273_t is
  variable rv : uint1273_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1273_t_to_slv(x : int1273_t) return std_logic_vector is
  variable rv : std_logic_vector(1272 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1273_t(x : std_logic_vector) return int1273_t is
  variable rv : int1273_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1274_t_to_slv(x : uint1274_t) return std_logic_vector is
  variable rv : std_logic_vector(1273 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1274_t(x : std_logic_vector) return uint1274_t is
  variable rv : uint1274_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1274_t_to_slv(x : int1274_t) return std_logic_vector is
  variable rv : std_logic_vector(1273 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1274_t(x : std_logic_vector) return int1274_t is
  variable rv : int1274_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1275_t_to_slv(x : uint1275_t) return std_logic_vector is
  variable rv : std_logic_vector(1274 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1275_t(x : std_logic_vector) return uint1275_t is
  variable rv : uint1275_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1275_t_to_slv(x : int1275_t) return std_logic_vector is
  variable rv : std_logic_vector(1274 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1275_t(x : std_logic_vector) return int1275_t is
  variable rv : int1275_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1276_t_to_slv(x : uint1276_t) return std_logic_vector is
  variable rv : std_logic_vector(1275 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1276_t(x : std_logic_vector) return uint1276_t is
  variable rv : uint1276_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1276_t_to_slv(x : int1276_t) return std_logic_vector is
  variable rv : std_logic_vector(1275 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1276_t(x : std_logic_vector) return int1276_t is
  variable rv : int1276_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1277_t_to_slv(x : uint1277_t) return std_logic_vector is
  variable rv : std_logic_vector(1276 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1277_t(x : std_logic_vector) return uint1277_t is
  variable rv : uint1277_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1277_t_to_slv(x : int1277_t) return std_logic_vector is
  variable rv : std_logic_vector(1276 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1277_t(x : std_logic_vector) return int1277_t is
  variable rv : int1277_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1278_t_to_slv(x : uint1278_t) return std_logic_vector is
  variable rv : std_logic_vector(1277 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1278_t(x : std_logic_vector) return uint1278_t is
  variable rv : uint1278_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1278_t_to_slv(x : int1278_t) return std_logic_vector is
  variable rv : std_logic_vector(1277 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1278_t(x : std_logic_vector) return int1278_t is
  variable rv : int1278_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1279_t_to_slv(x : uint1279_t) return std_logic_vector is
  variable rv : std_logic_vector(1278 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1279_t(x : std_logic_vector) return uint1279_t is
  variable rv : uint1279_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1279_t_to_slv(x : int1279_t) return std_logic_vector is
  variable rv : std_logic_vector(1278 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1279_t(x : std_logic_vector) return int1279_t is
  variable rv : int1279_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1280_t_to_slv(x : uint1280_t) return std_logic_vector is
  variable rv : std_logic_vector(1279 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1280_t(x : std_logic_vector) return uint1280_t is
  variable rv : uint1280_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1280_t_to_slv(x : int1280_t) return std_logic_vector is
  variable rv : std_logic_vector(1279 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1280_t(x : std_logic_vector) return int1280_t is
  variable rv : int1280_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1281_t_to_slv(x : uint1281_t) return std_logic_vector is
  variable rv : std_logic_vector(1280 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1281_t(x : std_logic_vector) return uint1281_t is
  variable rv : uint1281_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1281_t_to_slv(x : int1281_t) return std_logic_vector is
  variable rv : std_logic_vector(1280 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1281_t(x : std_logic_vector) return int1281_t is
  variable rv : int1281_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1282_t_to_slv(x : uint1282_t) return std_logic_vector is
  variable rv : std_logic_vector(1281 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1282_t(x : std_logic_vector) return uint1282_t is
  variable rv : uint1282_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1282_t_to_slv(x : int1282_t) return std_logic_vector is
  variable rv : std_logic_vector(1281 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1282_t(x : std_logic_vector) return int1282_t is
  variable rv : int1282_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1283_t_to_slv(x : uint1283_t) return std_logic_vector is
  variable rv : std_logic_vector(1282 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1283_t(x : std_logic_vector) return uint1283_t is
  variable rv : uint1283_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1283_t_to_slv(x : int1283_t) return std_logic_vector is
  variable rv : std_logic_vector(1282 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1283_t(x : std_logic_vector) return int1283_t is
  variable rv : int1283_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1284_t_to_slv(x : uint1284_t) return std_logic_vector is
  variable rv : std_logic_vector(1283 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1284_t(x : std_logic_vector) return uint1284_t is
  variable rv : uint1284_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1284_t_to_slv(x : int1284_t) return std_logic_vector is
  variable rv : std_logic_vector(1283 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1284_t(x : std_logic_vector) return int1284_t is
  variable rv : int1284_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1285_t_to_slv(x : uint1285_t) return std_logic_vector is
  variable rv : std_logic_vector(1284 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1285_t(x : std_logic_vector) return uint1285_t is
  variable rv : uint1285_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1285_t_to_slv(x : int1285_t) return std_logic_vector is
  variable rv : std_logic_vector(1284 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1285_t(x : std_logic_vector) return int1285_t is
  variable rv : int1285_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1286_t_to_slv(x : uint1286_t) return std_logic_vector is
  variable rv : std_logic_vector(1285 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1286_t(x : std_logic_vector) return uint1286_t is
  variable rv : uint1286_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1286_t_to_slv(x : int1286_t) return std_logic_vector is
  variable rv : std_logic_vector(1285 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1286_t(x : std_logic_vector) return int1286_t is
  variable rv : int1286_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1287_t_to_slv(x : uint1287_t) return std_logic_vector is
  variable rv : std_logic_vector(1286 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1287_t(x : std_logic_vector) return uint1287_t is
  variable rv : uint1287_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1287_t_to_slv(x : int1287_t) return std_logic_vector is
  variable rv : std_logic_vector(1286 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1287_t(x : std_logic_vector) return int1287_t is
  variable rv : int1287_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1288_t_to_slv(x : uint1288_t) return std_logic_vector is
  variable rv : std_logic_vector(1287 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1288_t(x : std_logic_vector) return uint1288_t is
  variable rv : uint1288_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1288_t_to_slv(x : int1288_t) return std_logic_vector is
  variable rv : std_logic_vector(1287 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1288_t(x : std_logic_vector) return int1288_t is
  variable rv : int1288_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1289_t_to_slv(x : uint1289_t) return std_logic_vector is
  variable rv : std_logic_vector(1288 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1289_t(x : std_logic_vector) return uint1289_t is
  variable rv : uint1289_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1289_t_to_slv(x : int1289_t) return std_logic_vector is
  variable rv : std_logic_vector(1288 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1289_t(x : std_logic_vector) return int1289_t is
  variable rv : int1289_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1290_t_to_slv(x : uint1290_t) return std_logic_vector is
  variable rv : std_logic_vector(1289 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1290_t(x : std_logic_vector) return uint1290_t is
  variable rv : uint1290_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1290_t_to_slv(x : int1290_t) return std_logic_vector is
  variable rv : std_logic_vector(1289 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1290_t(x : std_logic_vector) return int1290_t is
  variable rv : int1290_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1291_t_to_slv(x : uint1291_t) return std_logic_vector is
  variable rv : std_logic_vector(1290 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1291_t(x : std_logic_vector) return uint1291_t is
  variable rv : uint1291_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1291_t_to_slv(x : int1291_t) return std_logic_vector is
  variable rv : std_logic_vector(1290 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1291_t(x : std_logic_vector) return int1291_t is
  variable rv : int1291_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1292_t_to_slv(x : uint1292_t) return std_logic_vector is
  variable rv : std_logic_vector(1291 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1292_t(x : std_logic_vector) return uint1292_t is
  variable rv : uint1292_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1292_t_to_slv(x : int1292_t) return std_logic_vector is
  variable rv : std_logic_vector(1291 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1292_t(x : std_logic_vector) return int1292_t is
  variable rv : int1292_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1293_t_to_slv(x : uint1293_t) return std_logic_vector is
  variable rv : std_logic_vector(1292 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1293_t(x : std_logic_vector) return uint1293_t is
  variable rv : uint1293_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1293_t_to_slv(x : int1293_t) return std_logic_vector is
  variable rv : std_logic_vector(1292 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1293_t(x : std_logic_vector) return int1293_t is
  variable rv : int1293_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1294_t_to_slv(x : uint1294_t) return std_logic_vector is
  variable rv : std_logic_vector(1293 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1294_t(x : std_logic_vector) return uint1294_t is
  variable rv : uint1294_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1294_t_to_slv(x : int1294_t) return std_logic_vector is
  variable rv : std_logic_vector(1293 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1294_t(x : std_logic_vector) return int1294_t is
  variable rv : int1294_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1295_t_to_slv(x : uint1295_t) return std_logic_vector is
  variable rv : std_logic_vector(1294 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1295_t(x : std_logic_vector) return uint1295_t is
  variable rv : uint1295_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1295_t_to_slv(x : int1295_t) return std_logic_vector is
  variable rv : std_logic_vector(1294 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1295_t(x : std_logic_vector) return int1295_t is
  variable rv : int1295_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1296_t_to_slv(x : uint1296_t) return std_logic_vector is
  variable rv : std_logic_vector(1295 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1296_t(x : std_logic_vector) return uint1296_t is
  variable rv : uint1296_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1296_t_to_slv(x : int1296_t) return std_logic_vector is
  variable rv : std_logic_vector(1295 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1296_t(x : std_logic_vector) return int1296_t is
  variable rv : int1296_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1297_t_to_slv(x : uint1297_t) return std_logic_vector is
  variable rv : std_logic_vector(1296 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1297_t(x : std_logic_vector) return uint1297_t is
  variable rv : uint1297_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1297_t_to_slv(x : int1297_t) return std_logic_vector is
  variable rv : std_logic_vector(1296 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1297_t(x : std_logic_vector) return int1297_t is
  variable rv : int1297_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1298_t_to_slv(x : uint1298_t) return std_logic_vector is
  variable rv : std_logic_vector(1297 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1298_t(x : std_logic_vector) return uint1298_t is
  variable rv : uint1298_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1298_t_to_slv(x : int1298_t) return std_logic_vector is
  variable rv : std_logic_vector(1297 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1298_t(x : std_logic_vector) return int1298_t is
  variable rv : int1298_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1299_t_to_slv(x : uint1299_t) return std_logic_vector is
  variable rv : std_logic_vector(1298 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1299_t(x : std_logic_vector) return uint1299_t is
  variable rv : uint1299_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1299_t_to_slv(x : int1299_t) return std_logic_vector is
  variable rv : std_logic_vector(1298 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1299_t(x : std_logic_vector) return int1299_t is
  variable rv : int1299_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1300_t_to_slv(x : uint1300_t) return std_logic_vector is
  variable rv : std_logic_vector(1299 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1300_t(x : std_logic_vector) return uint1300_t is
  variable rv : uint1300_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1300_t_to_slv(x : int1300_t) return std_logic_vector is
  variable rv : std_logic_vector(1299 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1300_t(x : std_logic_vector) return int1300_t is
  variable rv : int1300_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1301_t_to_slv(x : uint1301_t) return std_logic_vector is
  variable rv : std_logic_vector(1300 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1301_t(x : std_logic_vector) return uint1301_t is
  variable rv : uint1301_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1301_t_to_slv(x : int1301_t) return std_logic_vector is
  variable rv : std_logic_vector(1300 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1301_t(x : std_logic_vector) return int1301_t is
  variable rv : int1301_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1302_t_to_slv(x : uint1302_t) return std_logic_vector is
  variable rv : std_logic_vector(1301 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1302_t(x : std_logic_vector) return uint1302_t is
  variable rv : uint1302_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1302_t_to_slv(x : int1302_t) return std_logic_vector is
  variable rv : std_logic_vector(1301 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1302_t(x : std_logic_vector) return int1302_t is
  variable rv : int1302_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1303_t_to_slv(x : uint1303_t) return std_logic_vector is
  variable rv : std_logic_vector(1302 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1303_t(x : std_logic_vector) return uint1303_t is
  variable rv : uint1303_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1303_t_to_slv(x : int1303_t) return std_logic_vector is
  variable rv : std_logic_vector(1302 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1303_t(x : std_logic_vector) return int1303_t is
  variable rv : int1303_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1304_t_to_slv(x : uint1304_t) return std_logic_vector is
  variable rv : std_logic_vector(1303 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1304_t(x : std_logic_vector) return uint1304_t is
  variable rv : uint1304_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1304_t_to_slv(x : int1304_t) return std_logic_vector is
  variable rv : std_logic_vector(1303 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1304_t(x : std_logic_vector) return int1304_t is
  variable rv : int1304_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1305_t_to_slv(x : uint1305_t) return std_logic_vector is
  variable rv : std_logic_vector(1304 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1305_t(x : std_logic_vector) return uint1305_t is
  variable rv : uint1305_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1305_t_to_slv(x : int1305_t) return std_logic_vector is
  variable rv : std_logic_vector(1304 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1305_t(x : std_logic_vector) return int1305_t is
  variable rv : int1305_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1306_t_to_slv(x : uint1306_t) return std_logic_vector is
  variable rv : std_logic_vector(1305 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1306_t(x : std_logic_vector) return uint1306_t is
  variable rv : uint1306_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1306_t_to_slv(x : int1306_t) return std_logic_vector is
  variable rv : std_logic_vector(1305 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1306_t(x : std_logic_vector) return int1306_t is
  variable rv : int1306_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1307_t_to_slv(x : uint1307_t) return std_logic_vector is
  variable rv : std_logic_vector(1306 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1307_t(x : std_logic_vector) return uint1307_t is
  variable rv : uint1307_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1307_t_to_slv(x : int1307_t) return std_logic_vector is
  variable rv : std_logic_vector(1306 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1307_t(x : std_logic_vector) return int1307_t is
  variable rv : int1307_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1308_t_to_slv(x : uint1308_t) return std_logic_vector is
  variable rv : std_logic_vector(1307 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1308_t(x : std_logic_vector) return uint1308_t is
  variable rv : uint1308_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1308_t_to_slv(x : int1308_t) return std_logic_vector is
  variable rv : std_logic_vector(1307 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1308_t(x : std_logic_vector) return int1308_t is
  variable rv : int1308_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1309_t_to_slv(x : uint1309_t) return std_logic_vector is
  variable rv : std_logic_vector(1308 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1309_t(x : std_logic_vector) return uint1309_t is
  variable rv : uint1309_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1309_t_to_slv(x : int1309_t) return std_logic_vector is
  variable rv : std_logic_vector(1308 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1309_t(x : std_logic_vector) return int1309_t is
  variable rv : int1309_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1310_t_to_slv(x : uint1310_t) return std_logic_vector is
  variable rv : std_logic_vector(1309 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1310_t(x : std_logic_vector) return uint1310_t is
  variable rv : uint1310_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1310_t_to_slv(x : int1310_t) return std_logic_vector is
  variable rv : std_logic_vector(1309 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1310_t(x : std_logic_vector) return int1310_t is
  variable rv : int1310_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1311_t_to_slv(x : uint1311_t) return std_logic_vector is
  variable rv : std_logic_vector(1310 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1311_t(x : std_logic_vector) return uint1311_t is
  variable rv : uint1311_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1311_t_to_slv(x : int1311_t) return std_logic_vector is
  variable rv : std_logic_vector(1310 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1311_t(x : std_logic_vector) return int1311_t is
  variable rv : int1311_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1312_t_to_slv(x : uint1312_t) return std_logic_vector is
  variable rv : std_logic_vector(1311 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1312_t(x : std_logic_vector) return uint1312_t is
  variable rv : uint1312_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1312_t_to_slv(x : int1312_t) return std_logic_vector is
  variable rv : std_logic_vector(1311 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1312_t(x : std_logic_vector) return int1312_t is
  variable rv : int1312_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1313_t_to_slv(x : uint1313_t) return std_logic_vector is
  variable rv : std_logic_vector(1312 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1313_t(x : std_logic_vector) return uint1313_t is
  variable rv : uint1313_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1313_t_to_slv(x : int1313_t) return std_logic_vector is
  variable rv : std_logic_vector(1312 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1313_t(x : std_logic_vector) return int1313_t is
  variable rv : int1313_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1314_t_to_slv(x : uint1314_t) return std_logic_vector is
  variable rv : std_logic_vector(1313 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1314_t(x : std_logic_vector) return uint1314_t is
  variable rv : uint1314_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1314_t_to_slv(x : int1314_t) return std_logic_vector is
  variable rv : std_logic_vector(1313 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1314_t(x : std_logic_vector) return int1314_t is
  variable rv : int1314_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1315_t_to_slv(x : uint1315_t) return std_logic_vector is
  variable rv : std_logic_vector(1314 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1315_t(x : std_logic_vector) return uint1315_t is
  variable rv : uint1315_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1315_t_to_slv(x : int1315_t) return std_logic_vector is
  variable rv : std_logic_vector(1314 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1315_t(x : std_logic_vector) return int1315_t is
  variable rv : int1315_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1316_t_to_slv(x : uint1316_t) return std_logic_vector is
  variable rv : std_logic_vector(1315 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1316_t(x : std_logic_vector) return uint1316_t is
  variable rv : uint1316_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1316_t_to_slv(x : int1316_t) return std_logic_vector is
  variable rv : std_logic_vector(1315 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1316_t(x : std_logic_vector) return int1316_t is
  variable rv : int1316_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1317_t_to_slv(x : uint1317_t) return std_logic_vector is
  variable rv : std_logic_vector(1316 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1317_t(x : std_logic_vector) return uint1317_t is
  variable rv : uint1317_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1317_t_to_slv(x : int1317_t) return std_logic_vector is
  variable rv : std_logic_vector(1316 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1317_t(x : std_logic_vector) return int1317_t is
  variable rv : int1317_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1318_t_to_slv(x : uint1318_t) return std_logic_vector is
  variable rv : std_logic_vector(1317 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1318_t(x : std_logic_vector) return uint1318_t is
  variable rv : uint1318_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1318_t_to_slv(x : int1318_t) return std_logic_vector is
  variable rv : std_logic_vector(1317 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1318_t(x : std_logic_vector) return int1318_t is
  variable rv : int1318_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1319_t_to_slv(x : uint1319_t) return std_logic_vector is
  variable rv : std_logic_vector(1318 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1319_t(x : std_logic_vector) return uint1319_t is
  variable rv : uint1319_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1319_t_to_slv(x : int1319_t) return std_logic_vector is
  variable rv : std_logic_vector(1318 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1319_t(x : std_logic_vector) return int1319_t is
  variable rv : int1319_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1320_t_to_slv(x : uint1320_t) return std_logic_vector is
  variable rv : std_logic_vector(1319 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1320_t(x : std_logic_vector) return uint1320_t is
  variable rv : uint1320_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1320_t_to_slv(x : int1320_t) return std_logic_vector is
  variable rv : std_logic_vector(1319 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1320_t(x : std_logic_vector) return int1320_t is
  variable rv : int1320_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1321_t_to_slv(x : uint1321_t) return std_logic_vector is
  variable rv : std_logic_vector(1320 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1321_t(x : std_logic_vector) return uint1321_t is
  variable rv : uint1321_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1321_t_to_slv(x : int1321_t) return std_logic_vector is
  variable rv : std_logic_vector(1320 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1321_t(x : std_logic_vector) return int1321_t is
  variable rv : int1321_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1322_t_to_slv(x : uint1322_t) return std_logic_vector is
  variable rv : std_logic_vector(1321 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1322_t(x : std_logic_vector) return uint1322_t is
  variable rv : uint1322_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1322_t_to_slv(x : int1322_t) return std_logic_vector is
  variable rv : std_logic_vector(1321 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1322_t(x : std_logic_vector) return int1322_t is
  variable rv : int1322_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1323_t_to_slv(x : uint1323_t) return std_logic_vector is
  variable rv : std_logic_vector(1322 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1323_t(x : std_logic_vector) return uint1323_t is
  variable rv : uint1323_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1323_t_to_slv(x : int1323_t) return std_logic_vector is
  variable rv : std_logic_vector(1322 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1323_t(x : std_logic_vector) return int1323_t is
  variable rv : int1323_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1324_t_to_slv(x : uint1324_t) return std_logic_vector is
  variable rv : std_logic_vector(1323 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1324_t(x : std_logic_vector) return uint1324_t is
  variable rv : uint1324_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1324_t_to_slv(x : int1324_t) return std_logic_vector is
  variable rv : std_logic_vector(1323 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1324_t(x : std_logic_vector) return int1324_t is
  variable rv : int1324_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1325_t_to_slv(x : uint1325_t) return std_logic_vector is
  variable rv : std_logic_vector(1324 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1325_t(x : std_logic_vector) return uint1325_t is
  variable rv : uint1325_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1325_t_to_slv(x : int1325_t) return std_logic_vector is
  variable rv : std_logic_vector(1324 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1325_t(x : std_logic_vector) return int1325_t is
  variable rv : int1325_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1326_t_to_slv(x : uint1326_t) return std_logic_vector is
  variable rv : std_logic_vector(1325 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1326_t(x : std_logic_vector) return uint1326_t is
  variable rv : uint1326_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1326_t_to_slv(x : int1326_t) return std_logic_vector is
  variable rv : std_logic_vector(1325 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1326_t(x : std_logic_vector) return int1326_t is
  variable rv : int1326_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1327_t_to_slv(x : uint1327_t) return std_logic_vector is
  variable rv : std_logic_vector(1326 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1327_t(x : std_logic_vector) return uint1327_t is
  variable rv : uint1327_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1327_t_to_slv(x : int1327_t) return std_logic_vector is
  variable rv : std_logic_vector(1326 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1327_t(x : std_logic_vector) return int1327_t is
  variable rv : int1327_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1328_t_to_slv(x : uint1328_t) return std_logic_vector is
  variable rv : std_logic_vector(1327 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1328_t(x : std_logic_vector) return uint1328_t is
  variable rv : uint1328_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1328_t_to_slv(x : int1328_t) return std_logic_vector is
  variable rv : std_logic_vector(1327 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1328_t(x : std_logic_vector) return int1328_t is
  variable rv : int1328_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1329_t_to_slv(x : uint1329_t) return std_logic_vector is
  variable rv : std_logic_vector(1328 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1329_t(x : std_logic_vector) return uint1329_t is
  variable rv : uint1329_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1329_t_to_slv(x : int1329_t) return std_logic_vector is
  variable rv : std_logic_vector(1328 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1329_t(x : std_logic_vector) return int1329_t is
  variable rv : int1329_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1330_t_to_slv(x : uint1330_t) return std_logic_vector is
  variable rv : std_logic_vector(1329 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1330_t(x : std_logic_vector) return uint1330_t is
  variable rv : uint1330_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1330_t_to_slv(x : int1330_t) return std_logic_vector is
  variable rv : std_logic_vector(1329 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1330_t(x : std_logic_vector) return int1330_t is
  variable rv : int1330_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1331_t_to_slv(x : uint1331_t) return std_logic_vector is
  variable rv : std_logic_vector(1330 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1331_t(x : std_logic_vector) return uint1331_t is
  variable rv : uint1331_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1331_t_to_slv(x : int1331_t) return std_logic_vector is
  variable rv : std_logic_vector(1330 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1331_t(x : std_logic_vector) return int1331_t is
  variable rv : int1331_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1332_t_to_slv(x : uint1332_t) return std_logic_vector is
  variable rv : std_logic_vector(1331 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1332_t(x : std_logic_vector) return uint1332_t is
  variable rv : uint1332_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1332_t_to_slv(x : int1332_t) return std_logic_vector is
  variable rv : std_logic_vector(1331 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1332_t(x : std_logic_vector) return int1332_t is
  variable rv : int1332_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1333_t_to_slv(x : uint1333_t) return std_logic_vector is
  variable rv : std_logic_vector(1332 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1333_t(x : std_logic_vector) return uint1333_t is
  variable rv : uint1333_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1333_t_to_slv(x : int1333_t) return std_logic_vector is
  variable rv : std_logic_vector(1332 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1333_t(x : std_logic_vector) return int1333_t is
  variable rv : int1333_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1334_t_to_slv(x : uint1334_t) return std_logic_vector is
  variable rv : std_logic_vector(1333 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1334_t(x : std_logic_vector) return uint1334_t is
  variable rv : uint1334_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1334_t_to_slv(x : int1334_t) return std_logic_vector is
  variable rv : std_logic_vector(1333 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1334_t(x : std_logic_vector) return int1334_t is
  variable rv : int1334_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1335_t_to_slv(x : uint1335_t) return std_logic_vector is
  variable rv : std_logic_vector(1334 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1335_t(x : std_logic_vector) return uint1335_t is
  variable rv : uint1335_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1335_t_to_slv(x : int1335_t) return std_logic_vector is
  variable rv : std_logic_vector(1334 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1335_t(x : std_logic_vector) return int1335_t is
  variable rv : int1335_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1336_t_to_slv(x : uint1336_t) return std_logic_vector is
  variable rv : std_logic_vector(1335 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1336_t(x : std_logic_vector) return uint1336_t is
  variable rv : uint1336_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1336_t_to_slv(x : int1336_t) return std_logic_vector is
  variable rv : std_logic_vector(1335 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1336_t(x : std_logic_vector) return int1336_t is
  variable rv : int1336_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1337_t_to_slv(x : uint1337_t) return std_logic_vector is
  variable rv : std_logic_vector(1336 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1337_t(x : std_logic_vector) return uint1337_t is
  variable rv : uint1337_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1337_t_to_slv(x : int1337_t) return std_logic_vector is
  variable rv : std_logic_vector(1336 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1337_t(x : std_logic_vector) return int1337_t is
  variable rv : int1337_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1338_t_to_slv(x : uint1338_t) return std_logic_vector is
  variable rv : std_logic_vector(1337 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1338_t(x : std_logic_vector) return uint1338_t is
  variable rv : uint1338_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1338_t_to_slv(x : int1338_t) return std_logic_vector is
  variable rv : std_logic_vector(1337 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1338_t(x : std_logic_vector) return int1338_t is
  variable rv : int1338_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1339_t_to_slv(x : uint1339_t) return std_logic_vector is
  variable rv : std_logic_vector(1338 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1339_t(x : std_logic_vector) return uint1339_t is
  variable rv : uint1339_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1339_t_to_slv(x : int1339_t) return std_logic_vector is
  variable rv : std_logic_vector(1338 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1339_t(x : std_logic_vector) return int1339_t is
  variable rv : int1339_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1340_t_to_slv(x : uint1340_t) return std_logic_vector is
  variable rv : std_logic_vector(1339 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1340_t(x : std_logic_vector) return uint1340_t is
  variable rv : uint1340_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1340_t_to_slv(x : int1340_t) return std_logic_vector is
  variable rv : std_logic_vector(1339 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1340_t(x : std_logic_vector) return int1340_t is
  variable rv : int1340_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1341_t_to_slv(x : uint1341_t) return std_logic_vector is
  variable rv : std_logic_vector(1340 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1341_t(x : std_logic_vector) return uint1341_t is
  variable rv : uint1341_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1341_t_to_slv(x : int1341_t) return std_logic_vector is
  variable rv : std_logic_vector(1340 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1341_t(x : std_logic_vector) return int1341_t is
  variable rv : int1341_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1342_t_to_slv(x : uint1342_t) return std_logic_vector is
  variable rv : std_logic_vector(1341 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1342_t(x : std_logic_vector) return uint1342_t is
  variable rv : uint1342_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1342_t_to_slv(x : int1342_t) return std_logic_vector is
  variable rv : std_logic_vector(1341 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1342_t(x : std_logic_vector) return int1342_t is
  variable rv : int1342_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1343_t_to_slv(x : uint1343_t) return std_logic_vector is
  variable rv : std_logic_vector(1342 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1343_t(x : std_logic_vector) return uint1343_t is
  variable rv : uint1343_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1343_t_to_slv(x : int1343_t) return std_logic_vector is
  variable rv : std_logic_vector(1342 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1343_t(x : std_logic_vector) return int1343_t is
  variable rv : int1343_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1344_t_to_slv(x : uint1344_t) return std_logic_vector is
  variable rv : std_logic_vector(1343 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1344_t(x : std_logic_vector) return uint1344_t is
  variable rv : uint1344_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1344_t_to_slv(x : int1344_t) return std_logic_vector is
  variable rv : std_logic_vector(1343 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1344_t(x : std_logic_vector) return int1344_t is
  variable rv : int1344_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1345_t_to_slv(x : uint1345_t) return std_logic_vector is
  variable rv : std_logic_vector(1344 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1345_t(x : std_logic_vector) return uint1345_t is
  variable rv : uint1345_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1345_t_to_slv(x : int1345_t) return std_logic_vector is
  variable rv : std_logic_vector(1344 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1345_t(x : std_logic_vector) return int1345_t is
  variable rv : int1345_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1346_t_to_slv(x : uint1346_t) return std_logic_vector is
  variable rv : std_logic_vector(1345 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1346_t(x : std_logic_vector) return uint1346_t is
  variable rv : uint1346_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1346_t_to_slv(x : int1346_t) return std_logic_vector is
  variable rv : std_logic_vector(1345 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1346_t(x : std_logic_vector) return int1346_t is
  variable rv : int1346_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1347_t_to_slv(x : uint1347_t) return std_logic_vector is
  variable rv : std_logic_vector(1346 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1347_t(x : std_logic_vector) return uint1347_t is
  variable rv : uint1347_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1347_t_to_slv(x : int1347_t) return std_logic_vector is
  variable rv : std_logic_vector(1346 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1347_t(x : std_logic_vector) return int1347_t is
  variable rv : int1347_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1348_t_to_slv(x : uint1348_t) return std_logic_vector is
  variable rv : std_logic_vector(1347 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1348_t(x : std_logic_vector) return uint1348_t is
  variable rv : uint1348_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1348_t_to_slv(x : int1348_t) return std_logic_vector is
  variable rv : std_logic_vector(1347 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1348_t(x : std_logic_vector) return int1348_t is
  variable rv : int1348_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1349_t_to_slv(x : uint1349_t) return std_logic_vector is
  variable rv : std_logic_vector(1348 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1349_t(x : std_logic_vector) return uint1349_t is
  variable rv : uint1349_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1349_t_to_slv(x : int1349_t) return std_logic_vector is
  variable rv : std_logic_vector(1348 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1349_t(x : std_logic_vector) return int1349_t is
  variable rv : int1349_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1350_t_to_slv(x : uint1350_t) return std_logic_vector is
  variable rv : std_logic_vector(1349 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1350_t(x : std_logic_vector) return uint1350_t is
  variable rv : uint1350_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1350_t_to_slv(x : int1350_t) return std_logic_vector is
  variable rv : std_logic_vector(1349 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1350_t(x : std_logic_vector) return int1350_t is
  variable rv : int1350_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1351_t_to_slv(x : uint1351_t) return std_logic_vector is
  variable rv : std_logic_vector(1350 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1351_t(x : std_logic_vector) return uint1351_t is
  variable rv : uint1351_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1351_t_to_slv(x : int1351_t) return std_logic_vector is
  variable rv : std_logic_vector(1350 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1351_t(x : std_logic_vector) return int1351_t is
  variable rv : int1351_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1352_t_to_slv(x : uint1352_t) return std_logic_vector is
  variable rv : std_logic_vector(1351 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1352_t(x : std_logic_vector) return uint1352_t is
  variable rv : uint1352_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1352_t_to_slv(x : int1352_t) return std_logic_vector is
  variable rv : std_logic_vector(1351 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1352_t(x : std_logic_vector) return int1352_t is
  variable rv : int1352_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1353_t_to_slv(x : uint1353_t) return std_logic_vector is
  variable rv : std_logic_vector(1352 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1353_t(x : std_logic_vector) return uint1353_t is
  variable rv : uint1353_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1353_t_to_slv(x : int1353_t) return std_logic_vector is
  variable rv : std_logic_vector(1352 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1353_t(x : std_logic_vector) return int1353_t is
  variable rv : int1353_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1354_t_to_slv(x : uint1354_t) return std_logic_vector is
  variable rv : std_logic_vector(1353 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1354_t(x : std_logic_vector) return uint1354_t is
  variable rv : uint1354_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1354_t_to_slv(x : int1354_t) return std_logic_vector is
  variable rv : std_logic_vector(1353 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1354_t(x : std_logic_vector) return int1354_t is
  variable rv : int1354_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1355_t_to_slv(x : uint1355_t) return std_logic_vector is
  variable rv : std_logic_vector(1354 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1355_t(x : std_logic_vector) return uint1355_t is
  variable rv : uint1355_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1355_t_to_slv(x : int1355_t) return std_logic_vector is
  variable rv : std_logic_vector(1354 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1355_t(x : std_logic_vector) return int1355_t is
  variable rv : int1355_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1356_t_to_slv(x : uint1356_t) return std_logic_vector is
  variable rv : std_logic_vector(1355 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1356_t(x : std_logic_vector) return uint1356_t is
  variable rv : uint1356_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1356_t_to_slv(x : int1356_t) return std_logic_vector is
  variable rv : std_logic_vector(1355 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1356_t(x : std_logic_vector) return int1356_t is
  variable rv : int1356_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1357_t_to_slv(x : uint1357_t) return std_logic_vector is
  variable rv : std_logic_vector(1356 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1357_t(x : std_logic_vector) return uint1357_t is
  variable rv : uint1357_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1357_t_to_slv(x : int1357_t) return std_logic_vector is
  variable rv : std_logic_vector(1356 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1357_t(x : std_logic_vector) return int1357_t is
  variable rv : int1357_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1358_t_to_slv(x : uint1358_t) return std_logic_vector is
  variable rv : std_logic_vector(1357 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1358_t(x : std_logic_vector) return uint1358_t is
  variable rv : uint1358_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1358_t_to_slv(x : int1358_t) return std_logic_vector is
  variable rv : std_logic_vector(1357 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1358_t(x : std_logic_vector) return int1358_t is
  variable rv : int1358_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1359_t_to_slv(x : uint1359_t) return std_logic_vector is
  variable rv : std_logic_vector(1358 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1359_t(x : std_logic_vector) return uint1359_t is
  variable rv : uint1359_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1359_t_to_slv(x : int1359_t) return std_logic_vector is
  variable rv : std_logic_vector(1358 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1359_t(x : std_logic_vector) return int1359_t is
  variable rv : int1359_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1360_t_to_slv(x : uint1360_t) return std_logic_vector is
  variable rv : std_logic_vector(1359 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1360_t(x : std_logic_vector) return uint1360_t is
  variable rv : uint1360_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1360_t_to_slv(x : int1360_t) return std_logic_vector is
  variable rv : std_logic_vector(1359 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1360_t(x : std_logic_vector) return int1360_t is
  variable rv : int1360_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1361_t_to_slv(x : uint1361_t) return std_logic_vector is
  variable rv : std_logic_vector(1360 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1361_t(x : std_logic_vector) return uint1361_t is
  variable rv : uint1361_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1361_t_to_slv(x : int1361_t) return std_logic_vector is
  variable rv : std_logic_vector(1360 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1361_t(x : std_logic_vector) return int1361_t is
  variable rv : int1361_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1362_t_to_slv(x : uint1362_t) return std_logic_vector is
  variable rv : std_logic_vector(1361 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1362_t(x : std_logic_vector) return uint1362_t is
  variable rv : uint1362_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1362_t_to_slv(x : int1362_t) return std_logic_vector is
  variable rv : std_logic_vector(1361 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1362_t(x : std_logic_vector) return int1362_t is
  variable rv : int1362_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1363_t_to_slv(x : uint1363_t) return std_logic_vector is
  variable rv : std_logic_vector(1362 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1363_t(x : std_logic_vector) return uint1363_t is
  variable rv : uint1363_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1363_t_to_slv(x : int1363_t) return std_logic_vector is
  variable rv : std_logic_vector(1362 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1363_t(x : std_logic_vector) return int1363_t is
  variable rv : int1363_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1364_t_to_slv(x : uint1364_t) return std_logic_vector is
  variable rv : std_logic_vector(1363 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1364_t(x : std_logic_vector) return uint1364_t is
  variable rv : uint1364_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1364_t_to_slv(x : int1364_t) return std_logic_vector is
  variable rv : std_logic_vector(1363 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1364_t(x : std_logic_vector) return int1364_t is
  variable rv : int1364_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1365_t_to_slv(x : uint1365_t) return std_logic_vector is
  variable rv : std_logic_vector(1364 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1365_t(x : std_logic_vector) return uint1365_t is
  variable rv : uint1365_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1365_t_to_slv(x : int1365_t) return std_logic_vector is
  variable rv : std_logic_vector(1364 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1365_t(x : std_logic_vector) return int1365_t is
  variable rv : int1365_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1366_t_to_slv(x : uint1366_t) return std_logic_vector is
  variable rv : std_logic_vector(1365 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1366_t(x : std_logic_vector) return uint1366_t is
  variable rv : uint1366_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1366_t_to_slv(x : int1366_t) return std_logic_vector is
  variable rv : std_logic_vector(1365 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1366_t(x : std_logic_vector) return int1366_t is
  variable rv : int1366_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1367_t_to_slv(x : uint1367_t) return std_logic_vector is
  variable rv : std_logic_vector(1366 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1367_t(x : std_logic_vector) return uint1367_t is
  variable rv : uint1367_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1367_t_to_slv(x : int1367_t) return std_logic_vector is
  variable rv : std_logic_vector(1366 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1367_t(x : std_logic_vector) return int1367_t is
  variable rv : int1367_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1368_t_to_slv(x : uint1368_t) return std_logic_vector is
  variable rv : std_logic_vector(1367 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1368_t(x : std_logic_vector) return uint1368_t is
  variable rv : uint1368_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1368_t_to_slv(x : int1368_t) return std_logic_vector is
  variable rv : std_logic_vector(1367 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1368_t(x : std_logic_vector) return int1368_t is
  variable rv : int1368_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1369_t_to_slv(x : uint1369_t) return std_logic_vector is
  variable rv : std_logic_vector(1368 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1369_t(x : std_logic_vector) return uint1369_t is
  variable rv : uint1369_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1369_t_to_slv(x : int1369_t) return std_logic_vector is
  variable rv : std_logic_vector(1368 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1369_t(x : std_logic_vector) return int1369_t is
  variable rv : int1369_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1370_t_to_slv(x : uint1370_t) return std_logic_vector is
  variable rv : std_logic_vector(1369 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1370_t(x : std_logic_vector) return uint1370_t is
  variable rv : uint1370_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1370_t_to_slv(x : int1370_t) return std_logic_vector is
  variable rv : std_logic_vector(1369 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1370_t(x : std_logic_vector) return int1370_t is
  variable rv : int1370_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1371_t_to_slv(x : uint1371_t) return std_logic_vector is
  variable rv : std_logic_vector(1370 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1371_t(x : std_logic_vector) return uint1371_t is
  variable rv : uint1371_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1371_t_to_slv(x : int1371_t) return std_logic_vector is
  variable rv : std_logic_vector(1370 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1371_t(x : std_logic_vector) return int1371_t is
  variable rv : int1371_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1372_t_to_slv(x : uint1372_t) return std_logic_vector is
  variable rv : std_logic_vector(1371 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1372_t(x : std_logic_vector) return uint1372_t is
  variable rv : uint1372_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1372_t_to_slv(x : int1372_t) return std_logic_vector is
  variable rv : std_logic_vector(1371 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1372_t(x : std_logic_vector) return int1372_t is
  variable rv : int1372_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1373_t_to_slv(x : uint1373_t) return std_logic_vector is
  variable rv : std_logic_vector(1372 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1373_t(x : std_logic_vector) return uint1373_t is
  variable rv : uint1373_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1373_t_to_slv(x : int1373_t) return std_logic_vector is
  variable rv : std_logic_vector(1372 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1373_t(x : std_logic_vector) return int1373_t is
  variable rv : int1373_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1374_t_to_slv(x : uint1374_t) return std_logic_vector is
  variable rv : std_logic_vector(1373 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1374_t(x : std_logic_vector) return uint1374_t is
  variable rv : uint1374_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1374_t_to_slv(x : int1374_t) return std_logic_vector is
  variable rv : std_logic_vector(1373 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1374_t(x : std_logic_vector) return int1374_t is
  variable rv : int1374_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1375_t_to_slv(x : uint1375_t) return std_logic_vector is
  variable rv : std_logic_vector(1374 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1375_t(x : std_logic_vector) return uint1375_t is
  variable rv : uint1375_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1375_t_to_slv(x : int1375_t) return std_logic_vector is
  variable rv : std_logic_vector(1374 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1375_t(x : std_logic_vector) return int1375_t is
  variable rv : int1375_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1376_t_to_slv(x : uint1376_t) return std_logic_vector is
  variable rv : std_logic_vector(1375 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1376_t(x : std_logic_vector) return uint1376_t is
  variable rv : uint1376_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1376_t_to_slv(x : int1376_t) return std_logic_vector is
  variable rv : std_logic_vector(1375 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1376_t(x : std_logic_vector) return int1376_t is
  variable rv : int1376_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1377_t_to_slv(x : uint1377_t) return std_logic_vector is
  variable rv : std_logic_vector(1376 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1377_t(x : std_logic_vector) return uint1377_t is
  variable rv : uint1377_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1377_t_to_slv(x : int1377_t) return std_logic_vector is
  variable rv : std_logic_vector(1376 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1377_t(x : std_logic_vector) return int1377_t is
  variable rv : int1377_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1378_t_to_slv(x : uint1378_t) return std_logic_vector is
  variable rv : std_logic_vector(1377 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1378_t(x : std_logic_vector) return uint1378_t is
  variable rv : uint1378_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1378_t_to_slv(x : int1378_t) return std_logic_vector is
  variable rv : std_logic_vector(1377 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1378_t(x : std_logic_vector) return int1378_t is
  variable rv : int1378_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1379_t_to_slv(x : uint1379_t) return std_logic_vector is
  variable rv : std_logic_vector(1378 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1379_t(x : std_logic_vector) return uint1379_t is
  variable rv : uint1379_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1379_t_to_slv(x : int1379_t) return std_logic_vector is
  variable rv : std_logic_vector(1378 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1379_t(x : std_logic_vector) return int1379_t is
  variable rv : int1379_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1380_t_to_slv(x : uint1380_t) return std_logic_vector is
  variable rv : std_logic_vector(1379 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1380_t(x : std_logic_vector) return uint1380_t is
  variable rv : uint1380_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1380_t_to_slv(x : int1380_t) return std_logic_vector is
  variable rv : std_logic_vector(1379 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1380_t(x : std_logic_vector) return int1380_t is
  variable rv : int1380_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1381_t_to_slv(x : uint1381_t) return std_logic_vector is
  variable rv : std_logic_vector(1380 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1381_t(x : std_logic_vector) return uint1381_t is
  variable rv : uint1381_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1381_t_to_slv(x : int1381_t) return std_logic_vector is
  variable rv : std_logic_vector(1380 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1381_t(x : std_logic_vector) return int1381_t is
  variable rv : int1381_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1382_t_to_slv(x : uint1382_t) return std_logic_vector is
  variable rv : std_logic_vector(1381 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1382_t(x : std_logic_vector) return uint1382_t is
  variable rv : uint1382_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1382_t_to_slv(x : int1382_t) return std_logic_vector is
  variable rv : std_logic_vector(1381 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1382_t(x : std_logic_vector) return int1382_t is
  variable rv : int1382_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1383_t_to_slv(x : uint1383_t) return std_logic_vector is
  variable rv : std_logic_vector(1382 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1383_t(x : std_logic_vector) return uint1383_t is
  variable rv : uint1383_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1383_t_to_slv(x : int1383_t) return std_logic_vector is
  variable rv : std_logic_vector(1382 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1383_t(x : std_logic_vector) return int1383_t is
  variable rv : int1383_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1384_t_to_slv(x : uint1384_t) return std_logic_vector is
  variable rv : std_logic_vector(1383 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1384_t(x : std_logic_vector) return uint1384_t is
  variable rv : uint1384_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1384_t_to_slv(x : int1384_t) return std_logic_vector is
  variable rv : std_logic_vector(1383 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1384_t(x : std_logic_vector) return int1384_t is
  variable rv : int1384_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1385_t_to_slv(x : uint1385_t) return std_logic_vector is
  variable rv : std_logic_vector(1384 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1385_t(x : std_logic_vector) return uint1385_t is
  variable rv : uint1385_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1385_t_to_slv(x : int1385_t) return std_logic_vector is
  variable rv : std_logic_vector(1384 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1385_t(x : std_logic_vector) return int1385_t is
  variable rv : int1385_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1386_t_to_slv(x : uint1386_t) return std_logic_vector is
  variable rv : std_logic_vector(1385 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1386_t(x : std_logic_vector) return uint1386_t is
  variable rv : uint1386_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1386_t_to_slv(x : int1386_t) return std_logic_vector is
  variable rv : std_logic_vector(1385 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1386_t(x : std_logic_vector) return int1386_t is
  variable rv : int1386_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1387_t_to_slv(x : uint1387_t) return std_logic_vector is
  variable rv : std_logic_vector(1386 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1387_t(x : std_logic_vector) return uint1387_t is
  variable rv : uint1387_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1387_t_to_slv(x : int1387_t) return std_logic_vector is
  variable rv : std_logic_vector(1386 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1387_t(x : std_logic_vector) return int1387_t is
  variable rv : int1387_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1388_t_to_slv(x : uint1388_t) return std_logic_vector is
  variable rv : std_logic_vector(1387 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1388_t(x : std_logic_vector) return uint1388_t is
  variable rv : uint1388_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1388_t_to_slv(x : int1388_t) return std_logic_vector is
  variable rv : std_logic_vector(1387 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1388_t(x : std_logic_vector) return int1388_t is
  variable rv : int1388_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1389_t_to_slv(x : uint1389_t) return std_logic_vector is
  variable rv : std_logic_vector(1388 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1389_t(x : std_logic_vector) return uint1389_t is
  variable rv : uint1389_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1389_t_to_slv(x : int1389_t) return std_logic_vector is
  variable rv : std_logic_vector(1388 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1389_t(x : std_logic_vector) return int1389_t is
  variable rv : int1389_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1390_t_to_slv(x : uint1390_t) return std_logic_vector is
  variable rv : std_logic_vector(1389 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1390_t(x : std_logic_vector) return uint1390_t is
  variable rv : uint1390_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1390_t_to_slv(x : int1390_t) return std_logic_vector is
  variable rv : std_logic_vector(1389 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1390_t(x : std_logic_vector) return int1390_t is
  variable rv : int1390_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1391_t_to_slv(x : uint1391_t) return std_logic_vector is
  variable rv : std_logic_vector(1390 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1391_t(x : std_logic_vector) return uint1391_t is
  variable rv : uint1391_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1391_t_to_slv(x : int1391_t) return std_logic_vector is
  variable rv : std_logic_vector(1390 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1391_t(x : std_logic_vector) return int1391_t is
  variable rv : int1391_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1392_t_to_slv(x : uint1392_t) return std_logic_vector is
  variable rv : std_logic_vector(1391 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1392_t(x : std_logic_vector) return uint1392_t is
  variable rv : uint1392_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1392_t_to_slv(x : int1392_t) return std_logic_vector is
  variable rv : std_logic_vector(1391 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1392_t(x : std_logic_vector) return int1392_t is
  variable rv : int1392_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1393_t_to_slv(x : uint1393_t) return std_logic_vector is
  variable rv : std_logic_vector(1392 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1393_t(x : std_logic_vector) return uint1393_t is
  variable rv : uint1393_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1393_t_to_slv(x : int1393_t) return std_logic_vector is
  variable rv : std_logic_vector(1392 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1393_t(x : std_logic_vector) return int1393_t is
  variable rv : int1393_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1394_t_to_slv(x : uint1394_t) return std_logic_vector is
  variable rv : std_logic_vector(1393 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1394_t(x : std_logic_vector) return uint1394_t is
  variable rv : uint1394_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1394_t_to_slv(x : int1394_t) return std_logic_vector is
  variable rv : std_logic_vector(1393 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1394_t(x : std_logic_vector) return int1394_t is
  variable rv : int1394_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1395_t_to_slv(x : uint1395_t) return std_logic_vector is
  variable rv : std_logic_vector(1394 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1395_t(x : std_logic_vector) return uint1395_t is
  variable rv : uint1395_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1395_t_to_slv(x : int1395_t) return std_logic_vector is
  variable rv : std_logic_vector(1394 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1395_t(x : std_logic_vector) return int1395_t is
  variable rv : int1395_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1396_t_to_slv(x : uint1396_t) return std_logic_vector is
  variable rv : std_logic_vector(1395 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1396_t(x : std_logic_vector) return uint1396_t is
  variable rv : uint1396_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1396_t_to_slv(x : int1396_t) return std_logic_vector is
  variable rv : std_logic_vector(1395 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1396_t(x : std_logic_vector) return int1396_t is
  variable rv : int1396_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1397_t_to_slv(x : uint1397_t) return std_logic_vector is
  variable rv : std_logic_vector(1396 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1397_t(x : std_logic_vector) return uint1397_t is
  variable rv : uint1397_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1397_t_to_slv(x : int1397_t) return std_logic_vector is
  variable rv : std_logic_vector(1396 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1397_t(x : std_logic_vector) return int1397_t is
  variable rv : int1397_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1398_t_to_slv(x : uint1398_t) return std_logic_vector is
  variable rv : std_logic_vector(1397 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1398_t(x : std_logic_vector) return uint1398_t is
  variable rv : uint1398_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1398_t_to_slv(x : int1398_t) return std_logic_vector is
  variable rv : std_logic_vector(1397 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1398_t(x : std_logic_vector) return int1398_t is
  variable rv : int1398_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1399_t_to_slv(x : uint1399_t) return std_logic_vector is
  variable rv : std_logic_vector(1398 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1399_t(x : std_logic_vector) return uint1399_t is
  variable rv : uint1399_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1399_t_to_slv(x : int1399_t) return std_logic_vector is
  variable rv : std_logic_vector(1398 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1399_t(x : std_logic_vector) return int1399_t is
  variable rv : int1399_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1400_t_to_slv(x : uint1400_t) return std_logic_vector is
  variable rv : std_logic_vector(1399 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1400_t(x : std_logic_vector) return uint1400_t is
  variable rv : uint1400_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1400_t_to_slv(x : int1400_t) return std_logic_vector is
  variable rv : std_logic_vector(1399 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1400_t(x : std_logic_vector) return int1400_t is
  variable rv : int1400_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1401_t_to_slv(x : uint1401_t) return std_logic_vector is
  variable rv : std_logic_vector(1400 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1401_t(x : std_logic_vector) return uint1401_t is
  variable rv : uint1401_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1401_t_to_slv(x : int1401_t) return std_logic_vector is
  variable rv : std_logic_vector(1400 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1401_t(x : std_logic_vector) return int1401_t is
  variable rv : int1401_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1402_t_to_slv(x : uint1402_t) return std_logic_vector is
  variable rv : std_logic_vector(1401 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1402_t(x : std_logic_vector) return uint1402_t is
  variable rv : uint1402_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1402_t_to_slv(x : int1402_t) return std_logic_vector is
  variable rv : std_logic_vector(1401 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1402_t(x : std_logic_vector) return int1402_t is
  variable rv : int1402_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1403_t_to_slv(x : uint1403_t) return std_logic_vector is
  variable rv : std_logic_vector(1402 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1403_t(x : std_logic_vector) return uint1403_t is
  variable rv : uint1403_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1403_t_to_slv(x : int1403_t) return std_logic_vector is
  variable rv : std_logic_vector(1402 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1403_t(x : std_logic_vector) return int1403_t is
  variable rv : int1403_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1404_t_to_slv(x : uint1404_t) return std_logic_vector is
  variable rv : std_logic_vector(1403 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1404_t(x : std_logic_vector) return uint1404_t is
  variable rv : uint1404_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1404_t_to_slv(x : int1404_t) return std_logic_vector is
  variable rv : std_logic_vector(1403 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1404_t(x : std_logic_vector) return int1404_t is
  variable rv : int1404_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1405_t_to_slv(x : uint1405_t) return std_logic_vector is
  variable rv : std_logic_vector(1404 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1405_t(x : std_logic_vector) return uint1405_t is
  variable rv : uint1405_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1405_t_to_slv(x : int1405_t) return std_logic_vector is
  variable rv : std_logic_vector(1404 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1405_t(x : std_logic_vector) return int1405_t is
  variable rv : int1405_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1406_t_to_slv(x : uint1406_t) return std_logic_vector is
  variable rv : std_logic_vector(1405 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1406_t(x : std_logic_vector) return uint1406_t is
  variable rv : uint1406_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1406_t_to_slv(x : int1406_t) return std_logic_vector is
  variable rv : std_logic_vector(1405 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1406_t(x : std_logic_vector) return int1406_t is
  variable rv : int1406_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1407_t_to_slv(x : uint1407_t) return std_logic_vector is
  variable rv : std_logic_vector(1406 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1407_t(x : std_logic_vector) return uint1407_t is
  variable rv : uint1407_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1407_t_to_slv(x : int1407_t) return std_logic_vector is
  variable rv : std_logic_vector(1406 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1407_t(x : std_logic_vector) return int1407_t is
  variable rv : int1407_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1408_t_to_slv(x : uint1408_t) return std_logic_vector is
  variable rv : std_logic_vector(1407 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1408_t(x : std_logic_vector) return uint1408_t is
  variable rv : uint1408_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1408_t_to_slv(x : int1408_t) return std_logic_vector is
  variable rv : std_logic_vector(1407 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1408_t(x : std_logic_vector) return int1408_t is
  variable rv : int1408_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1409_t_to_slv(x : uint1409_t) return std_logic_vector is
  variable rv : std_logic_vector(1408 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1409_t(x : std_logic_vector) return uint1409_t is
  variable rv : uint1409_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1409_t_to_slv(x : int1409_t) return std_logic_vector is
  variable rv : std_logic_vector(1408 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1409_t(x : std_logic_vector) return int1409_t is
  variable rv : int1409_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1410_t_to_slv(x : uint1410_t) return std_logic_vector is
  variable rv : std_logic_vector(1409 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1410_t(x : std_logic_vector) return uint1410_t is
  variable rv : uint1410_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1410_t_to_slv(x : int1410_t) return std_logic_vector is
  variable rv : std_logic_vector(1409 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1410_t(x : std_logic_vector) return int1410_t is
  variable rv : int1410_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1411_t_to_slv(x : uint1411_t) return std_logic_vector is
  variable rv : std_logic_vector(1410 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1411_t(x : std_logic_vector) return uint1411_t is
  variable rv : uint1411_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1411_t_to_slv(x : int1411_t) return std_logic_vector is
  variable rv : std_logic_vector(1410 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1411_t(x : std_logic_vector) return int1411_t is
  variable rv : int1411_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1412_t_to_slv(x : uint1412_t) return std_logic_vector is
  variable rv : std_logic_vector(1411 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1412_t(x : std_logic_vector) return uint1412_t is
  variable rv : uint1412_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1412_t_to_slv(x : int1412_t) return std_logic_vector is
  variable rv : std_logic_vector(1411 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1412_t(x : std_logic_vector) return int1412_t is
  variable rv : int1412_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1413_t_to_slv(x : uint1413_t) return std_logic_vector is
  variable rv : std_logic_vector(1412 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1413_t(x : std_logic_vector) return uint1413_t is
  variable rv : uint1413_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1413_t_to_slv(x : int1413_t) return std_logic_vector is
  variable rv : std_logic_vector(1412 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1413_t(x : std_logic_vector) return int1413_t is
  variable rv : int1413_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1414_t_to_slv(x : uint1414_t) return std_logic_vector is
  variable rv : std_logic_vector(1413 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1414_t(x : std_logic_vector) return uint1414_t is
  variable rv : uint1414_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1414_t_to_slv(x : int1414_t) return std_logic_vector is
  variable rv : std_logic_vector(1413 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1414_t(x : std_logic_vector) return int1414_t is
  variable rv : int1414_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1415_t_to_slv(x : uint1415_t) return std_logic_vector is
  variable rv : std_logic_vector(1414 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1415_t(x : std_logic_vector) return uint1415_t is
  variable rv : uint1415_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1415_t_to_slv(x : int1415_t) return std_logic_vector is
  variable rv : std_logic_vector(1414 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1415_t(x : std_logic_vector) return int1415_t is
  variable rv : int1415_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1416_t_to_slv(x : uint1416_t) return std_logic_vector is
  variable rv : std_logic_vector(1415 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1416_t(x : std_logic_vector) return uint1416_t is
  variable rv : uint1416_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1416_t_to_slv(x : int1416_t) return std_logic_vector is
  variable rv : std_logic_vector(1415 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1416_t(x : std_logic_vector) return int1416_t is
  variable rv : int1416_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1417_t_to_slv(x : uint1417_t) return std_logic_vector is
  variable rv : std_logic_vector(1416 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1417_t(x : std_logic_vector) return uint1417_t is
  variable rv : uint1417_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1417_t_to_slv(x : int1417_t) return std_logic_vector is
  variable rv : std_logic_vector(1416 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1417_t(x : std_logic_vector) return int1417_t is
  variable rv : int1417_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1418_t_to_slv(x : uint1418_t) return std_logic_vector is
  variable rv : std_logic_vector(1417 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1418_t(x : std_logic_vector) return uint1418_t is
  variable rv : uint1418_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1418_t_to_slv(x : int1418_t) return std_logic_vector is
  variable rv : std_logic_vector(1417 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1418_t(x : std_logic_vector) return int1418_t is
  variable rv : int1418_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1419_t_to_slv(x : uint1419_t) return std_logic_vector is
  variable rv : std_logic_vector(1418 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1419_t(x : std_logic_vector) return uint1419_t is
  variable rv : uint1419_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1419_t_to_slv(x : int1419_t) return std_logic_vector is
  variable rv : std_logic_vector(1418 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1419_t(x : std_logic_vector) return int1419_t is
  variable rv : int1419_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1420_t_to_slv(x : uint1420_t) return std_logic_vector is
  variable rv : std_logic_vector(1419 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1420_t(x : std_logic_vector) return uint1420_t is
  variable rv : uint1420_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1420_t_to_slv(x : int1420_t) return std_logic_vector is
  variable rv : std_logic_vector(1419 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1420_t(x : std_logic_vector) return int1420_t is
  variable rv : int1420_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1421_t_to_slv(x : uint1421_t) return std_logic_vector is
  variable rv : std_logic_vector(1420 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1421_t(x : std_logic_vector) return uint1421_t is
  variable rv : uint1421_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1421_t_to_slv(x : int1421_t) return std_logic_vector is
  variable rv : std_logic_vector(1420 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1421_t(x : std_logic_vector) return int1421_t is
  variable rv : int1421_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1422_t_to_slv(x : uint1422_t) return std_logic_vector is
  variable rv : std_logic_vector(1421 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1422_t(x : std_logic_vector) return uint1422_t is
  variable rv : uint1422_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1422_t_to_slv(x : int1422_t) return std_logic_vector is
  variable rv : std_logic_vector(1421 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1422_t(x : std_logic_vector) return int1422_t is
  variable rv : int1422_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1423_t_to_slv(x : uint1423_t) return std_logic_vector is
  variable rv : std_logic_vector(1422 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1423_t(x : std_logic_vector) return uint1423_t is
  variable rv : uint1423_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1423_t_to_slv(x : int1423_t) return std_logic_vector is
  variable rv : std_logic_vector(1422 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1423_t(x : std_logic_vector) return int1423_t is
  variable rv : int1423_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1424_t_to_slv(x : uint1424_t) return std_logic_vector is
  variable rv : std_logic_vector(1423 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1424_t(x : std_logic_vector) return uint1424_t is
  variable rv : uint1424_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1424_t_to_slv(x : int1424_t) return std_logic_vector is
  variable rv : std_logic_vector(1423 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1424_t(x : std_logic_vector) return int1424_t is
  variable rv : int1424_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1425_t_to_slv(x : uint1425_t) return std_logic_vector is
  variable rv : std_logic_vector(1424 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1425_t(x : std_logic_vector) return uint1425_t is
  variable rv : uint1425_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1425_t_to_slv(x : int1425_t) return std_logic_vector is
  variable rv : std_logic_vector(1424 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1425_t(x : std_logic_vector) return int1425_t is
  variable rv : int1425_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1426_t_to_slv(x : uint1426_t) return std_logic_vector is
  variable rv : std_logic_vector(1425 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1426_t(x : std_logic_vector) return uint1426_t is
  variable rv : uint1426_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1426_t_to_slv(x : int1426_t) return std_logic_vector is
  variable rv : std_logic_vector(1425 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1426_t(x : std_logic_vector) return int1426_t is
  variable rv : int1426_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1427_t_to_slv(x : uint1427_t) return std_logic_vector is
  variable rv : std_logic_vector(1426 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1427_t(x : std_logic_vector) return uint1427_t is
  variable rv : uint1427_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1427_t_to_slv(x : int1427_t) return std_logic_vector is
  variable rv : std_logic_vector(1426 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1427_t(x : std_logic_vector) return int1427_t is
  variable rv : int1427_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1428_t_to_slv(x : uint1428_t) return std_logic_vector is
  variable rv : std_logic_vector(1427 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1428_t(x : std_logic_vector) return uint1428_t is
  variable rv : uint1428_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1428_t_to_slv(x : int1428_t) return std_logic_vector is
  variable rv : std_logic_vector(1427 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1428_t(x : std_logic_vector) return int1428_t is
  variable rv : int1428_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1429_t_to_slv(x : uint1429_t) return std_logic_vector is
  variable rv : std_logic_vector(1428 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1429_t(x : std_logic_vector) return uint1429_t is
  variable rv : uint1429_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1429_t_to_slv(x : int1429_t) return std_logic_vector is
  variable rv : std_logic_vector(1428 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1429_t(x : std_logic_vector) return int1429_t is
  variable rv : int1429_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1430_t_to_slv(x : uint1430_t) return std_logic_vector is
  variable rv : std_logic_vector(1429 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1430_t(x : std_logic_vector) return uint1430_t is
  variable rv : uint1430_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1430_t_to_slv(x : int1430_t) return std_logic_vector is
  variable rv : std_logic_vector(1429 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1430_t(x : std_logic_vector) return int1430_t is
  variable rv : int1430_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1431_t_to_slv(x : uint1431_t) return std_logic_vector is
  variable rv : std_logic_vector(1430 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1431_t(x : std_logic_vector) return uint1431_t is
  variable rv : uint1431_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1431_t_to_slv(x : int1431_t) return std_logic_vector is
  variable rv : std_logic_vector(1430 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1431_t(x : std_logic_vector) return int1431_t is
  variable rv : int1431_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1432_t_to_slv(x : uint1432_t) return std_logic_vector is
  variable rv : std_logic_vector(1431 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1432_t(x : std_logic_vector) return uint1432_t is
  variable rv : uint1432_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1432_t_to_slv(x : int1432_t) return std_logic_vector is
  variable rv : std_logic_vector(1431 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1432_t(x : std_logic_vector) return int1432_t is
  variable rv : int1432_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1433_t_to_slv(x : uint1433_t) return std_logic_vector is
  variable rv : std_logic_vector(1432 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1433_t(x : std_logic_vector) return uint1433_t is
  variable rv : uint1433_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1433_t_to_slv(x : int1433_t) return std_logic_vector is
  variable rv : std_logic_vector(1432 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1433_t(x : std_logic_vector) return int1433_t is
  variable rv : int1433_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1434_t_to_slv(x : uint1434_t) return std_logic_vector is
  variable rv : std_logic_vector(1433 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1434_t(x : std_logic_vector) return uint1434_t is
  variable rv : uint1434_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1434_t_to_slv(x : int1434_t) return std_logic_vector is
  variable rv : std_logic_vector(1433 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1434_t(x : std_logic_vector) return int1434_t is
  variable rv : int1434_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1435_t_to_slv(x : uint1435_t) return std_logic_vector is
  variable rv : std_logic_vector(1434 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1435_t(x : std_logic_vector) return uint1435_t is
  variable rv : uint1435_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1435_t_to_slv(x : int1435_t) return std_logic_vector is
  variable rv : std_logic_vector(1434 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1435_t(x : std_logic_vector) return int1435_t is
  variable rv : int1435_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1436_t_to_slv(x : uint1436_t) return std_logic_vector is
  variable rv : std_logic_vector(1435 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1436_t(x : std_logic_vector) return uint1436_t is
  variable rv : uint1436_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1436_t_to_slv(x : int1436_t) return std_logic_vector is
  variable rv : std_logic_vector(1435 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1436_t(x : std_logic_vector) return int1436_t is
  variable rv : int1436_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1437_t_to_slv(x : uint1437_t) return std_logic_vector is
  variable rv : std_logic_vector(1436 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1437_t(x : std_logic_vector) return uint1437_t is
  variable rv : uint1437_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1437_t_to_slv(x : int1437_t) return std_logic_vector is
  variable rv : std_logic_vector(1436 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1437_t(x : std_logic_vector) return int1437_t is
  variable rv : int1437_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1438_t_to_slv(x : uint1438_t) return std_logic_vector is
  variable rv : std_logic_vector(1437 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1438_t(x : std_logic_vector) return uint1438_t is
  variable rv : uint1438_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1438_t_to_slv(x : int1438_t) return std_logic_vector is
  variable rv : std_logic_vector(1437 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1438_t(x : std_logic_vector) return int1438_t is
  variable rv : int1438_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1439_t_to_slv(x : uint1439_t) return std_logic_vector is
  variable rv : std_logic_vector(1438 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1439_t(x : std_logic_vector) return uint1439_t is
  variable rv : uint1439_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1439_t_to_slv(x : int1439_t) return std_logic_vector is
  variable rv : std_logic_vector(1438 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1439_t(x : std_logic_vector) return int1439_t is
  variable rv : int1439_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1440_t_to_slv(x : uint1440_t) return std_logic_vector is
  variable rv : std_logic_vector(1439 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1440_t(x : std_logic_vector) return uint1440_t is
  variable rv : uint1440_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1440_t_to_slv(x : int1440_t) return std_logic_vector is
  variable rv : std_logic_vector(1439 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1440_t(x : std_logic_vector) return int1440_t is
  variable rv : int1440_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1441_t_to_slv(x : uint1441_t) return std_logic_vector is
  variable rv : std_logic_vector(1440 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1441_t(x : std_logic_vector) return uint1441_t is
  variable rv : uint1441_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1441_t_to_slv(x : int1441_t) return std_logic_vector is
  variable rv : std_logic_vector(1440 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1441_t(x : std_logic_vector) return int1441_t is
  variable rv : int1441_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1442_t_to_slv(x : uint1442_t) return std_logic_vector is
  variable rv : std_logic_vector(1441 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1442_t(x : std_logic_vector) return uint1442_t is
  variable rv : uint1442_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1442_t_to_slv(x : int1442_t) return std_logic_vector is
  variable rv : std_logic_vector(1441 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1442_t(x : std_logic_vector) return int1442_t is
  variable rv : int1442_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1443_t_to_slv(x : uint1443_t) return std_logic_vector is
  variable rv : std_logic_vector(1442 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1443_t(x : std_logic_vector) return uint1443_t is
  variable rv : uint1443_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1443_t_to_slv(x : int1443_t) return std_logic_vector is
  variable rv : std_logic_vector(1442 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1443_t(x : std_logic_vector) return int1443_t is
  variable rv : int1443_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1444_t_to_slv(x : uint1444_t) return std_logic_vector is
  variable rv : std_logic_vector(1443 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1444_t(x : std_logic_vector) return uint1444_t is
  variable rv : uint1444_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1444_t_to_slv(x : int1444_t) return std_logic_vector is
  variable rv : std_logic_vector(1443 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1444_t(x : std_logic_vector) return int1444_t is
  variable rv : int1444_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1445_t_to_slv(x : uint1445_t) return std_logic_vector is
  variable rv : std_logic_vector(1444 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1445_t(x : std_logic_vector) return uint1445_t is
  variable rv : uint1445_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1445_t_to_slv(x : int1445_t) return std_logic_vector is
  variable rv : std_logic_vector(1444 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1445_t(x : std_logic_vector) return int1445_t is
  variable rv : int1445_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1446_t_to_slv(x : uint1446_t) return std_logic_vector is
  variable rv : std_logic_vector(1445 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1446_t(x : std_logic_vector) return uint1446_t is
  variable rv : uint1446_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1446_t_to_slv(x : int1446_t) return std_logic_vector is
  variable rv : std_logic_vector(1445 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1446_t(x : std_logic_vector) return int1446_t is
  variable rv : int1446_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1447_t_to_slv(x : uint1447_t) return std_logic_vector is
  variable rv : std_logic_vector(1446 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1447_t(x : std_logic_vector) return uint1447_t is
  variable rv : uint1447_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1447_t_to_slv(x : int1447_t) return std_logic_vector is
  variable rv : std_logic_vector(1446 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1447_t(x : std_logic_vector) return int1447_t is
  variable rv : int1447_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1448_t_to_slv(x : uint1448_t) return std_logic_vector is
  variable rv : std_logic_vector(1447 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1448_t(x : std_logic_vector) return uint1448_t is
  variable rv : uint1448_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1448_t_to_slv(x : int1448_t) return std_logic_vector is
  variable rv : std_logic_vector(1447 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1448_t(x : std_logic_vector) return int1448_t is
  variable rv : int1448_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1449_t_to_slv(x : uint1449_t) return std_logic_vector is
  variable rv : std_logic_vector(1448 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1449_t(x : std_logic_vector) return uint1449_t is
  variable rv : uint1449_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1449_t_to_slv(x : int1449_t) return std_logic_vector is
  variable rv : std_logic_vector(1448 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1449_t(x : std_logic_vector) return int1449_t is
  variable rv : int1449_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1450_t_to_slv(x : uint1450_t) return std_logic_vector is
  variable rv : std_logic_vector(1449 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1450_t(x : std_logic_vector) return uint1450_t is
  variable rv : uint1450_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1450_t_to_slv(x : int1450_t) return std_logic_vector is
  variable rv : std_logic_vector(1449 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1450_t(x : std_logic_vector) return int1450_t is
  variable rv : int1450_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1451_t_to_slv(x : uint1451_t) return std_logic_vector is
  variable rv : std_logic_vector(1450 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1451_t(x : std_logic_vector) return uint1451_t is
  variable rv : uint1451_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1451_t_to_slv(x : int1451_t) return std_logic_vector is
  variable rv : std_logic_vector(1450 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1451_t(x : std_logic_vector) return int1451_t is
  variable rv : int1451_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1452_t_to_slv(x : uint1452_t) return std_logic_vector is
  variable rv : std_logic_vector(1451 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1452_t(x : std_logic_vector) return uint1452_t is
  variable rv : uint1452_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1452_t_to_slv(x : int1452_t) return std_logic_vector is
  variable rv : std_logic_vector(1451 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1452_t(x : std_logic_vector) return int1452_t is
  variable rv : int1452_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1453_t_to_slv(x : uint1453_t) return std_logic_vector is
  variable rv : std_logic_vector(1452 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1453_t(x : std_logic_vector) return uint1453_t is
  variable rv : uint1453_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1453_t_to_slv(x : int1453_t) return std_logic_vector is
  variable rv : std_logic_vector(1452 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1453_t(x : std_logic_vector) return int1453_t is
  variable rv : int1453_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1454_t_to_slv(x : uint1454_t) return std_logic_vector is
  variable rv : std_logic_vector(1453 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1454_t(x : std_logic_vector) return uint1454_t is
  variable rv : uint1454_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1454_t_to_slv(x : int1454_t) return std_logic_vector is
  variable rv : std_logic_vector(1453 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1454_t(x : std_logic_vector) return int1454_t is
  variable rv : int1454_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1455_t_to_slv(x : uint1455_t) return std_logic_vector is
  variable rv : std_logic_vector(1454 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1455_t(x : std_logic_vector) return uint1455_t is
  variable rv : uint1455_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1455_t_to_slv(x : int1455_t) return std_logic_vector is
  variable rv : std_logic_vector(1454 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1455_t(x : std_logic_vector) return int1455_t is
  variable rv : int1455_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1456_t_to_slv(x : uint1456_t) return std_logic_vector is
  variable rv : std_logic_vector(1455 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1456_t(x : std_logic_vector) return uint1456_t is
  variable rv : uint1456_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1456_t_to_slv(x : int1456_t) return std_logic_vector is
  variable rv : std_logic_vector(1455 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1456_t(x : std_logic_vector) return int1456_t is
  variable rv : int1456_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1457_t_to_slv(x : uint1457_t) return std_logic_vector is
  variable rv : std_logic_vector(1456 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1457_t(x : std_logic_vector) return uint1457_t is
  variable rv : uint1457_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1457_t_to_slv(x : int1457_t) return std_logic_vector is
  variable rv : std_logic_vector(1456 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1457_t(x : std_logic_vector) return int1457_t is
  variable rv : int1457_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1458_t_to_slv(x : uint1458_t) return std_logic_vector is
  variable rv : std_logic_vector(1457 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1458_t(x : std_logic_vector) return uint1458_t is
  variable rv : uint1458_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1458_t_to_slv(x : int1458_t) return std_logic_vector is
  variable rv : std_logic_vector(1457 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1458_t(x : std_logic_vector) return int1458_t is
  variable rv : int1458_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1459_t_to_slv(x : uint1459_t) return std_logic_vector is
  variable rv : std_logic_vector(1458 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1459_t(x : std_logic_vector) return uint1459_t is
  variable rv : uint1459_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1459_t_to_slv(x : int1459_t) return std_logic_vector is
  variable rv : std_logic_vector(1458 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1459_t(x : std_logic_vector) return int1459_t is
  variable rv : int1459_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1460_t_to_slv(x : uint1460_t) return std_logic_vector is
  variable rv : std_logic_vector(1459 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1460_t(x : std_logic_vector) return uint1460_t is
  variable rv : uint1460_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1460_t_to_slv(x : int1460_t) return std_logic_vector is
  variable rv : std_logic_vector(1459 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1460_t(x : std_logic_vector) return int1460_t is
  variable rv : int1460_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1461_t_to_slv(x : uint1461_t) return std_logic_vector is
  variable rv : std_logic_vector(1460 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1461_t(x : std_logic_vector) return uint1461_t is
  variable rv : uint1461_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1461_t_to_slv(x : int1461_t) return std_logic_vector is
  variable rv : std_logic_vector(1460 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1461_t(x : std_logic_vector) return int1461_t is
  variable rv : int1461_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1462_t_to_slv(x : uint1462_t) return std_logic_vector is
  variable rv : std_logic_vector(1461 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1462_t(x : std_logic_vector) return uint1462_t is
  variable rv : uint1462_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1462_t_to_slv(x : int1462_t) return std_logic_vector is
  variable rv : std_logic_vector(1461 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1462_t(x : std_logic_vector) return int1462_t is
  variable rv : int1462_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1463_t_to_slv(x : uint1463_t) return std_logic_vector is
  variable rv : std_logic_vector(1462 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1463_t(x : std_logic_vector) return uint1463_t is
  variable rv : uint1463_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1463_t_to_slv(x : int1463_t) return std_logic_vector is
  variable rv : std_logic_vector(1462 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1463_t(x : std_logic_vector) return int1463_t is
  variable rv : int1463_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1464_t_to_slv(x : uint1464_t) return std_logic_vector is
  variable rv : std_logic_vector(1463 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1464_t(x : std_logic_vector) return uint1464_t is
  variable rv : uint1464_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1464_t_to_slv(x : int1464_t) return std_logic_vector is
  variable rv : std_logic_vector(1463 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1464_t(x : std_logic_vector) return int1464_t is
  variable rv : int1464_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1465_t_to_slv(x : uint1465_t) return std_logic_vector is
  variable rv : std_logic_vector(1464 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1465_t(x : std_logic_vector) return uint1465_t is
  variable rv : uint1465_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1465_t_to_slv(x : int1465_t) return std_logic_vector is
  variable rv : std_logic_vector(1464 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1465_t(x : std_logic_vector) return int1465_t is
  variable rv : int1465_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1466_t_to_slv(x : uint1466_t) return std_logic_vector is
  variable rv : std_logic_vector(1465 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1466_t(x : std_logic_vector) return uint1466_t is
  variable rv : uint1466_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1466_t_to_slv(x : int1466_t) return std_logic_vector is
  variable rv : std_logic_vector(1465 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1466_t(x : std_logic_vector) return int1466_t is
  variable rv : int1466_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1467_t_to_slv(x : uint1467_t) return std_logic_vector is
  variable rv : std_logic_vector(1466 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1467_t(x : std_logic_vector) return uint1467_t is
  variable rv : uint1467_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1467_t_to_slv(x : int1467_t) return std_logic_vector is
  variable rv : std_logic_vector(1466 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1467_t(x : std_logic_vector) return int1467_t is
  variable rv : int1467_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1468_t_to_slv(x : uint1468_t) return std_logic_vector is
  variable rv : std_logic_vector(1467 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1468_t(x : std_logic_vector) return uint1468_t is
  variable rv : uint1468_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1468_t_to_slv(x : int1468_t) return std_logic_vector is
  variable rv : std_logic_vector(1467 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1468_t(x : std_logic_vector) return int1468_t is
  variable rv : int1468_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1469_t_to_slv(x : uint1469_t) return std_logic_vector is
  variable rv : std_logic_vector(1468 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1469_t(x : std_logic_vector) return uint1469_t is
  variable rv : uint1469_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1469_t_to_slv(x : int1469_t) return std_logic_vector is
  variable rv : std_logic_vector(1468 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1469_t(x : std_logic_vector) return int1469_t is
  variable rv : int1469_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1470_t_to_slv(x : uint1470_t) return std_logic_vector is
  variable rv : std_logic_vector(1469 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1470_t(x : std_logic_vector) return uint1470_t is
  variable rv : uint1470_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1470_t_to_slv(x : int1470_t) return std_logic_vector is
  variable rv : std_logic_vector(1469 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1470_t(x : std_logic_vector) return int1470_t is
  variable rv : int1470_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1471_t_to_slv(x : uint1471_t) return std_logic_vector is
  variable rv : std_logic_vector(1470 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1471_t(x : std_logic_vector) return uint1471_t is
  variable rv : uint1471_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1471_t_to_slv(x : int1471_t) return std_logic_vector is
  variable rv : std_logic_vector(1470 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1471_t(x : std_logic_vector) return int1471_t is
  variable rv : int1471_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1472_t_to_slv(x : uint1472_t) return std_logic_vector is
  variable rv : std_logic_vector(1471 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1472_t(x : std_logic_vector) return uint1472_t is
  variable rv : uint1472_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1472_t_to_slv(x : int1472_t) return std_logic_vector is
  variable rv : std_logic_vector(1471 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1472_t(x : std_logic_vector) return int1472_t is
  variable rv : int1472_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1473_t_to_slv(x : uint1473_t) return std_logic_vector is
  variable rv : std_logic_vector(1472 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1473_t(x : std_logic_vector) return uint1473_t is
  variable rv : uint1473_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1473_t_to_slv(x : int1473_t) return std_logic_vector is
  variable rv : std_logic_vector(1472 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1473_t(x : std_logic_vector) return int1473_t is
  variable rv : int1473_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1474_t_to_slv(x : uint1474_t) return std_logic_vector is
  variable rv : std_logic_vector(1473 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1474_t(x : std_logic_vector) return uint1474_t is
  variable rv : uint1474_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1474_t_to_slv(x : int1474_t) return std_logic_vector is
  variable rv : std_logic_vector(1473 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1474_t(x : std_logic_vector) return int1474_t is
  variable rv : int1474_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1475_t_to_slv(x : uint1475_t) return std_logic_vector is
  variable rv : std_logic_vector(1474 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1475_t(x : std_logic_vector) return uint1475_t is
  variable rv : uint1475_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1475_t_to_slv(x : int1475_t) return std_logic_vector is
  variable rv : std_logic_vector(1474 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1475_t(x : std_logic_vector) return int1475_t is
  variable rv : int1475_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1476_t_to_slv(x : uint1476_t) return std_logic_vector is
  variable rv : std_logic_vector(1475 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1476_t(x : std_logic_vector) return uint1476_t is
  variable rv : uint1476_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1476_t_to_slv(x : int1476_t) return std_logic_vector is
  variable rv : std_logic_vector(1475 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1476_t(x : std_logic_vector) return int1476_t is
  variable rv : int1476_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1477_t_to_slv(x : uint1477_t) return std_logic_vector is
  variable rv : std_logic_vector(1476 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1477_t(x : std_logic_vector) return uint1477_t is
  variable rv : uint1477_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1477_t_to_slv(x : int1477_t) return std_logic_vector is
  variable rv : std_logic_vector(1476 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1477_t(x : std_logic_vector) return int1477_t is
  variable rv : int1477_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1478_t_to_slv(x : uint1478_t) return std_logic_vector is
  variable rv : std_logic_vector(1477 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1478_t(x : std_logic_vector) return uint1478_t is
  variable rv : uint1478_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1478_t_to_slv(x : int1478_t) return std_logic_vector is
  variable rv : std_logic_vector(1477 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1478_t(x : std_logic_vector) return int1478_t is
  variable rv : int1478_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1479_t_to_slv(x : uint1479_t) return std_logic_vector is
  variable rv : std_logic_vector(1478 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1479_t(x : std_logic_vector) return uint1479_t is
  variable rv : uint1479_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1479_t_to_slv(x : int1479_t) return std_logic_vector is
  variable rv : std_logic_vector(1478 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1479_t(x : std_logic_vector) return int1479_t is
  variable rv : int1479_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1480_t_to_slv(x : uint1480_t) return std_logic_vector is
  variable rv : std_logic_vector(1479 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1480_t(x : std_logic_vector) return uint1480_t is
  variable rv : uint1480_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1480_t_to_slv(x : int1480_t) return std_logic_vector is
  variable rv : std_logic_vector(1479 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1480_t(x : std_logic_vector) return int1480_t is
  variable rv : int1480_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1481_t_to_slv(x : uint1481_t) return std_logic_vector is
  variable rv : std_logic_vector(1480 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1481_t(x : std_logic_vector) return uint1481_t is
  variable rv : uint1481_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1481_t_to_slv(x : int1481_t) return std_logic_vector is
  variable rv : std_logic_vector(1480 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1481_t(x : std_logic_vector) return int1481_t is
  variable rv : int1481_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1482_t_to_slv(x : uint1482_t) return std_logic_vector is
  variable rv : std_logic_vector(1481 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1482_t(x : std_logic_vector) return uint1482_t is
  variable rv : uint1482_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1482_t_to_slv(x : int1482_t) return std_logic_vector is
  variable rv : std_logic_vector(1481 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1482_t(x : std_logic_vector) return int1482_t is
  variable rv : int1482_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1483_t_to_slv(x : uint1483_t) return std_logic_vector is
  variable rv : std_logic_vector(1482 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1483_t(x : std_logic_vector) return uint1483_t is
  variable rv : uint1483_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1483_t_to_slv(x : int1483_t) return std_logic_vector is
  variable rv : std_logic_vector(1482 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1483_t(x : std_logic_vector) return int1483_t is
  variable rv : int1483_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1484_t_to_slv(x : uint1484_t) return std_logic_vector is
  variable rv : std_logic_vector(1483 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1484_t(x : std_logic_vector) return uint1484_t is
  variable rv : uint1484_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1484_t_to_slv(x : int1484_t) return std_logic_vector is
  variable rv : std_logic_vector(1483 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1484_t(x : std_logic_vector) return int1484_t is
  variable rv : int1484_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1485_t_to_slv(x : uint1485_t) return std_logic_vector is
  variable rv : std_logic_vector(1484 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1485_t(x : std_logic_vector) return uint1485_t is
  variable rv : uint1485_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1485_t_to_slv(x : int1485_t) return std_logic_vector is
  variable rv : std_logic_vector(1484 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1485_t(x : std_logic_vector) return int1485_t is
  variable rv : int1485_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1486_t_to_slv(x : uint1486_t) return std_logic_vector is
  variable rv : std_logic_vector(1485 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1486_t(x : std_logic_vector) return uint1486_t is
  variable rv : uint1486_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1486_t_to_slv(x : int1486_t) return std_logic_vector is
  variable rv : std_logic_vector(1485 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1486_t(x : std_logic_vector) return int1486_t is
  variable rv : int1486_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1487_t_to_slv(x : uint1487_t) return std_logic_vector is
  variable rv : std_logic_vector(1486 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1487_t(x : std_logic_vector) return uint1487_t is
  variable rv : uint1487_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1487_t_to_slv(x : int1487_t) return std_logic_vector is
  variable rv : std_logic_vector(1486 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1487_t(x : std_logic_vector) return int1487_t is
  variable rv : int1487_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1488_t_to_slv(x : uint1488_t) return std_logic_vector is
  variable rv : std_logic_vector(1487 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1488_t(x : std_logic_vector) return uint1488_t is
  variable rv : uint1488_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1488_t_to_slv(x : int1488_t) return std_logic_vector is
  variable rv : std_logic_vector(1487 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1488_t(x : std_logic_vector) return int1488_t is
  variable rv : int1488_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1489_t_to_slv(x : uint1489_t) return std_logic_vector is
  variable rv : std_logic_vector(1488 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1489_t(x : std_logic_vector) return uint1489_t is
  variable rv : uint1489_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1489_t_to_slv(x : int1489_t) return std_logic_vector is
  variable rv : std_logic_vector(1488 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1489_t(x : std_logic_vector) return int1489_t is
  variable rv : int1489_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1490_t_to_slv(x : uint1490_t) return std_logic_vector is
  variable rv : std_logic_vector(1489 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1490_t(x : std_logic_vector) return uint1490_t is
  variable rv : uint1490_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1490_t_to_slv(x : int1490_t) return std_logic_vector is
  variable rv : std_logic_vector(1489 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1490_t(x : std_logic_vector) return int1490_t is
  variable rv : int1490_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1491_t_to_slv(x : uint1491_t) return std_logic_vector is
  variable rv : std_logic_vector(1490 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1491_t(x : std_logic_vector) return uint1491_t is
  variable rv : uint1491_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1491_t_to_slv(x : int1491_t) return std_logic_vector is
  variable rv : std_logic_vector(1490 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1491_t(x : std_logic_vector) return int1491_t is
  variable rv : int1491_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1492_t_to_slv(x : uint1492_t) return std_logic_vector is
  variable rv : std_logic_vector(1491 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1492_t(x : std_logic_vector) return uint1492_t is
  variable rv : uint1492_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1492_t_to_slv(x : int1492_t) return std_logic_vector is
  variable rv : std_logic_vector(1491 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1492_t(x : std_logic_vector) return int1492_t is
  variable rv : int1492_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1493_t_to_slv(x : uint1493_t) return std_logic_vector is
  variable rv : std_logic_vector(1492 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1493_t(x : std_logic_vector) return uint1493_t is
  variable rv : uint1493_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1493_t_to_slv(x : int1493_t) return std_logic_vector is
  variable rv : std_logic_vector(1492 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1493_t(x : std_logic_vector) return int1493_t is
  variable rv : int1493_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1494_t_to_slv(x : uint1494_t) return std_logic_vector is
  variable rv : std_logic_vector(1493 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1494_t(x : std_logic_vector) return uint1494_t is
  variable rv : uint1494_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1494_t_to_slv(x : int1494_t) return std_logic_vector is
  variable rv : std_logic_vector(1493 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1494_t(x : std_logic_vector) return int1494_t is
  variable rv : int1494_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1495_t_to_slv(x : uint1495_t) return std_logic_vector is
  variable rv : std_logic_vector(1494 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1495_t(x : std_logic_vector) return uint1495_t is
  variable rv : uint1495_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1495_t_to_slv(x : int1495_t) return std_logic_vector is
  variable rv : std_logic_vector(1494 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1495_t(x : std_logic_vector) return int1495_t is
  variable rv : int1495_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1496_t_to_slv(x : uint1496_t) return std_logic_vector is
  variable rv : std_logic_vector(1495 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1496_t(x : std_logic_vector) return uint1496_t is
  variable rv : uint1496_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1496_t_to_slv(x : int1496_t) return std_logic_vector is
  variable rv : std_logic_vector(1495 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1496_t(x : std_logic_vector) return int1496_t is
  variable rv : int1496_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1497_t_to_slv(x : uint1497_t) return std_logic_vector is
  variable rv : std_logic_vector(1496 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1497_t(x : std_logic_vector) return uint1497_t is
  variable rv : uint1497_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1497_t_to_slv(x : int1497_t) return std_logic_vector is
  variable rv : std_logic_vector(1496 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1497_t(x : std_logic_vector) return int1497_t is
  variable rv : int1497_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1498_t_to_slv(x : uint1498_t) return std_logic_vector is
  variable rv : std_logic_vector(1497 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1498_t(x : std_logic_vector) return uint1498_t is
  variable rv : uint1498_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1498_t_to_slv(x : int1498_t) return std_logic_vector is
  variable rv : std_logic_vector(1497 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1498_t(x : std_logic_vector) return int1498_t is
  variable rv : int1498_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1499_t_to_slv(x : uint1499_t) return std_logic_vector is
  variable rv : std_logic_vector(1498 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1499_t(x : std_logic_vector) return uint1499_t is
  variable rv : uint1499_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1499_t_to_slv(x : int1499_t) return std_logic_vector is
  variable rv : std_logic_vector(1498 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1499_t(x : std_logic_vector) return int1499_t is
  variable rv : int1499_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1500_t_to_slv(x : uint1500_t) return std_logic_vector is
  variable rv : std_logic_vector(1499 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1500_t(x : std_logic_vector) return uint1500_t is
  variable rv : uint1500_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1500_t_to_slv(x : int1500_t) return std_logic_vector is
  variable rv : std_logic_vector(1499 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1500_t(x : std_logic_vector) return int1500_t is
  variable rv : int1500_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1501_t_to_slv(x : uint1501_t) return std_logic_vector is
  variable rv : std_logic_vector(1500 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1501_t(x : std_logic_vector) return uint1501_t is
  variable rv : uint1501_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1501_t_to_slv(x : int1501_t) return std_logic_vector is
  variable rv : std_logic_vector(1500 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1501_t(x : std_logic_vector) return int1501_t is
  variable rv : int1501_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1502_t_to_slv(x : uint1502_t) return std_logic_vector is
  variable rv : std_logic_vector(1501 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1502_t(x : std_logic_vector) return uint1502_t is
  variable rv : uint1502_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1502_t_to_slv(x : int1502_t) return std_logic_vector is
  variable rv : std_logic_vector(1501 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1502_t(x : std_logic_vector) return int1502_t is
  variable rv : int1502_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1503_t_to_slv(x : uint1503_t) return std_logic_vector is
  variable rv : std_logic_vector(1502 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1503_t(x : std_logic_vector) return uint1503_t is
  variable rv : uint1503_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1503_t_to_slv(x : int1503_t) return std_logic_vector is
  variable rv : std_logic_vector(1502 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1503_t(x : std_logic_vector) return int1503_t is
  variable rv : int1503_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1504_t_to_slv(x : uint1504_t) return std_logic_vector is
  variable rv : std_logic_vector(1503 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1504_t(x : std_logic_vector) return uint1504_t is
  variable rv : uint1504_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1504_t_to_slv(x : int1504_t) return std_logic_vector is
  variable rv : std_logic_vector(1503 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1504_t(x : std_logic_vector) return int1504_t is
  variable rv : int1504_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1505_t_to_slv(x : uint1505_t) return std_logic_vector is
  variable rv : std_logic_vector(1504 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1505_t(x : std_logic_vector) return uint1505_t is
  variable rv : uint1505_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1505_t_to_slv(x : int1505_t) return std_logic_vector is
  variable rv : std_logic_vector(1504 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1505_t(x : std_logic_vector) return int1505_t is
  variable rv : int1505_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1506_t_to_slv(x : uint1506_t) return std_logic_vector is
  variable rv : std_logic_vector(1505 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1506_t(x : std_logic_vector) return uint1506_t is
  variable rv : uint1506_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1506_t_to_slv(x : int1506_t) return std_logic_vector is
  variable rv : std_logic_vector(1505 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1506_t(x : std_logic_vector) return int1506_t is
  variable rv : int1506_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1507_t_to_slv(x : uint1507_t) return std_logic_vector is
  variable rv : std_logic_vector(1506 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1507_t(x : std_logic_vector) return uint1507_t is
  variable rv : uint1507_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1507_t_to_slv(x : int1507_t) return std_logic_vector is
  variable rv : std_logic_vector(1506 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1507_t(x : std_logic_vector) return int1507_t is
  variable rv : int1507_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1508_t_to_slv(x : uint1508_t) return std_logic_vector is
  variable rv : std_logic_vector(1507 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1508_t(x : std_logic_vector) return uint1508_t is
  variable rv : uint1508_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1508_t_to_slv(x : int1508_t) return std_logic_vector is
  variable rv : std_logic_vector(1507 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1508_t(x : std_logic_vector) return int1508_t is
  variable rv : int1508_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1509_t_to_slv(x : uint1509_t) return std_logic_vector is
  variable rv : std_logic_vector(1508 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1509_t(x : std_logic_vector) return uint1509_t is
  variable rv : uint1509_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1509_t_to_slv(x : int1509_t) return std_logic_vector is
  variable rv : std_logic_vector(1508 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1509_t(x : std_logic_vector) return int1509_t is
  variable rv : int1509_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1510_t_to_slv(x : uint1510_t) return std_logic_vector is
  variable rv : std_logic_vector(1509 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1510_t(x : std_logic_vector) return uint1510_t is
  variable rv : uint1510_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1510_t_to_slv(x : int1510_t) return std_logic_vector is
  variable rv : std_logic_vector(1509 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1510_t(x : std_logic_vector) return int1510_t is
  variable rv : int1510_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1511_t_to_slv(x : uint1511_t) return std_logic_vector is
  variable rv : std_logic_vector(1510 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1511_t(x : std_logic_vector) return uint1511_t is
  variable rv : uint1511_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1511_t_to_slv(x : int1511_t) return std_logic_vector is
  variable rv : std_logic_vector(1510 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1511_t(x : std_logic_vector) return int1511_t is
  variable rv : int1511_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1512_t_to_slv(x : uint1512_t) return std_logic_vector is
  variable rv : std_logic_vector(1511 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1512_t(x : std_logic_vector) return uint1512_t is
  variable rv : uint1512_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1512_t_to_slv(x : int1512_t) return std_logic_vector is
  variable rv : std_logic_vector(1511 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1512_t(x : std_logic_vector) return int1512_t is
  variable rv : int1512_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1513_t_to_slv(x : uint1513_t) return std_logic_vector is
  variable rv : std_logic_vector(1512 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1513_t(x : std_logic_vector) return uint1513_t is
  variable rv : uint1513_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1513_t_to_slv(x : int1513_t) return std_logic_vector is
  variable rv : std_logic_vector(1512 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1513_t(x : std_logic_vector) return int1513_t is
  variable rv : int1513_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1514_t_to_slv(x : uint1514_t) return std_logic_vector is
  variable rv : std_logic_vector(1513 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1514_t(x : std_logic_vector) return uint1514_t is
  variable rv : uint1514_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1514_t_to_slv(x : int1514_t) return std_logic_vector is
  variable rv : std_logic_vector(1513 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1514_t(x : std_logic_vector) return int1514_t is
  variable rv : int1514_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1515_t_to_slv(x : uint1515_t) return std_logic_vector is
  variable rv : std_logic_vector(1514 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1515_t(x : std_logic_vector) return uint1515_t is
  variable rv : uint1515_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1515_t_to_slv(x : int1515_t) return std_logic_vector is
  variable rv : std_logic_vector(1514 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1515_t(x : std_logic_vector) return int1515_t is
  variable rv : int1515_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1516_t_to_slv(x : uint1516_t) return std_logic_vector is
  variable rv : std_logic_vector(1515 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1516_t(x : std_logic_vector) return uint1516_t is
  variable rv : uint1516_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1516_t_to_slv(x : int1516_t) return std_logic_vector is
  variable rv : std_logic_vector(1515 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1516_t(x : std_logic_vector) return int1516_t is
  variable rv : int1516_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1517_t_to_slv(x : uint1517_t) return std_logic_vector is
  variable rv : std_logic_vector(1516 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1517_t(x : std_logic_vector) return uint1517_t is
  variable rv : uint1517_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1517_t_to_slv(x : int1517_t) return std_logic_vector is
  variable rv : std_logic_vector(1516 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1517_t(x : std_logic_vector) return int1517_t is
  variable rv : int1517_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1518_t_to_slv(x : uint1518_t) return std_logic_vector is
  variable rv : std_logic_vector(1517 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1518_t(x : std_logic_vector) return uint1518_t is
  variable rv : uint1518_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1518_t_to_slv(x : int1518_t) return std_logic_vector is
  variable rv : std_logic_vector(1517 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1518_t(x : std_logic_vector) return int1518_t is
  variable rv : int1518_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1519_t_to_slv(x : uint1519_t) return std_logic_vector is
  variable rv : std_logic_vector(1518 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1519_t(x : std_logic_vector) return uint1519_t is
  variable rv : uint1519_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1519_t_to_slv(x : int1519_t) return std_logic_vector is
  variable rv : std_logic_vector(1518 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1519_t(x : std_logic_vector) return int1519_t is
  variable rv : int1519_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1520_t_to_slv(x : uint1520_t) return std_logic_vector is
  variable rv : std_logic_vector(1519 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1520_t(x : std_logic_vector) return uint1520_t is
  variable rv : uint1520_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1520_t_to_slv(x : int1520_t) return std_logic_vector is
  variable rv : std_logic_vector(1519 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1520_t(x : std_logic_vector) return int1520_t is
  variable rv : int1520_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1521_t_to_slv(x : uint1521_t) return std_logic_vector is
  variable rv : std_logic_vector(1520 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1521_t(x : std_logic_vector) return uint1521_t is
  variable rv : uint1521_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1521_t_to_slv(x : int1521_t) return std_logic_vector is
  variable rv : std_logic_vector(1520 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1521_t(x : std_logic_vector) return int1521_t is
  variable rv : int1521_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1522_t_to_slv(x : uint1522_t) return std_logic_vector is
  variable rv : std_logic_vector(1521 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1522_t(x : std_logic_vector) return uint1522_t is
  variable rv : uint1522_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1522_t_to_slv(x : int1522_t) return std_logic_vector is
  variable rv : std_logic_vector(1521 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1522_t(x : std_logic_vector) return int1522_t is
  variable rv : int1522_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1523_t_to_slv(x : uint1523_t) return std_logic_vector is
  variable rv : std_logic_vector(1522 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1523_t(x : std_logic_vector) return uint1523_t is
  variable rv : uint1523_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1523_t_to_slv(x : int1523_t) return std_logic_vector is
  variable rv : std_logic_vector(1522 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1523_t(x : std_logic_vector) return int1523_t is
  variable rv : int1523_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1524_t_to_slv(x : uint1524_t) return std_logic_vector is
  variable rv : std_logic_vector(1523 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1524_t(x : std_logic_vector) return uint1524_t is
  variable rv : uint1524_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1524_t_to_slv(x : int1524_t) return std_logic_vector is
  variable rv : std_logic_vector(1523 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1524_t(x : std_logic_vector) return int1524_t is
  variable rv : int1524_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1525_t_to_slv(x : uint1525_t) return std_logic_vector is
  variable rv : std_logic_vector(1524 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1525_t(x : std_logic_vector) return uint1525_t is
  variable rv : uint1525_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1525_t_to_slv(x : int1525_t) return std_logic_vector is
  variable rv : std_logic_vector(1524 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1525_t(x : std_logic_vector) return int1525_t is
  variable rv : int1525_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1526_t_to_slv(x : uint1526_t) return std_logic_vector is
  variable rv : std_logic_vector(1525 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1526_t(x : std_logic_vector) return uint1526_t is
  variable rv : uint1526_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1526_t_to_slv(x : int1526_t) return std_logic_vector is
  variable rv : std_logic_vector(1525 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1526_t(x : std_logic_vector) return int1526_t is
  variable rv : int1526_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1527_t_to_slv(x : uint1527_t) return std_logic_vector is
  variable rv : std_logic_vector(1526 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1527_t(x : std_logic_vector) return uint1527_t is
  variable rv : uint1527_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1527_t_to_slv(x : int1527_t) return std_logic_vector is
  variable rv : std_logic_vector(1526 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1527_t(x : std_logic_vector) return int1527_t is
  variable rv : int1527_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1528_t_to_slv(x : uint1528_t) return std_logic_vector is
  variable rv : std_logic_vector(1527 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1528_t(x : std_logic_vector) return uint1528_t is
  variable rv : uint1528_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1528_t_to_slv(x : int1528_t) return std_logic_vector is
  variable rv : std_logic_vector(1527 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1528_t(x : std_logic_vector) return int1528_t is
  variable rv : int1528_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1529_t_to_slv(x : uint1529_t) return std_logic_vector is
  variable rv : std_logic_vector(1528 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1529_t(x : std_logic_vector) return uint1529_t is
  variable rv : uint1529_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1529_t_to_slv(x : int1529_t) return std_logic_vector is
  variable rv : std_logic_vector(1528 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1529_t(x : std_logic_vector) return int1529_t is
  variable rv : int1529_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1530_t_to_slv(x : uint1530_t) return std_logic_vector is
  variable rv : std_logic_vector(1529 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1530_t(x : std_logic_vector) return uint1530_t is
  variable rv : uint1530_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1530_t_to_slv(x : int1530_t) return std_logic_vector is
  variable rv : std_logic_vector(1529 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1530_t(x : std_logic_vector) return int1530_t is
  variable rv : int1530_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1531_t_to_slv(x : uint1531_t) return std_logic_vector is
  variable rv : std_logic_vector(1530 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1531_t(x : std_logic_vector) return uint1531_t is
  variable rv : uint1531_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1531_t_to_slv(x : int1531_t) return std_logic_vector is
  variable rv : std_logic_vector(1530 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1531_t(x : std_logic_vector) return int1531_t is
  variable rv : int1531_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1532_t_to_slv(x : uint1532_t) return std_logic_vector is
  variable rv : std_logic_vector(1531 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1532_t(x : std_logic_vector) return uint1532_t is
  variable rv : uint1532_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1532_t_to_slv(x : int1532_t) return std_logic_vector is
  variable rv : std_logic_vector(1531 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1532_t(x : std_logic_vector) return int1532_t is
  variable rv : int1532_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1533_t_to_slv(x : uint1533_t) return std_logic_vector is
  variable rv : std_logic_vector(1532 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1533_t(x : std_logic_vector) return uint1533_t is
  variable rv : uint1533_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1533_t_to_slv(x : int1533_t) return std_logic_vector is
  variable rv : std_logic_vector(1532 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1533_t(x : std_logic_vector) return int1533_t is
  variable rv : int1533_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1534_t_to_slv(x : uint1534_t) return std_logic_vector is
  variable rv : std_logic_vector(1533 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1534_t(x : std_logic_vector) return uint1534_t is
  variable rv : uint1534_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1534_t_to_slv(x : int1534_t) return std_logic_vector is
  variable rv : std_logic_vector(1533 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1534_t(x : std_logic_vector) return int1534_t is
  variable rv : int1534_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1535_t_to_slv(x : uint1535_t) return std_logic_vector is
  variable rv : std_logic_vector(1534 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1535_t(x : std_logic_vector) return uint1535_t is
  variable rv : uint1535_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1535_t_to_slv(x : int1535_t) return std_logic_vector is
  variable rv : std_logic_vector(1534 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1535_t(x : std_logic_vector) return int1535_t is
  variable rv : int1535_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1536_t_to_slv(x : uint1536_t) return std_logic_vector is
  variable rv : std_logic_vector(1535 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1536_t(x : std_logic_vector) return uint1536_t is
  variable rv : uint1536_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1536_t_to_slv(x : int1536_t) return std_logic_vector is
  variable rv : std_logic_vector(1535 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1536_t(x : std_logic_vector) return int1536_t is
  variable rv : int1536_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1537_t_to_slv(x : uint1537_t) return std_logic_vector is
  variable rv : std_logic_vector(1536 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1537_t(x : std_logic_vector) return uint1537_t is
  variable rv : uint1537_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1537_t_to_slv(x : int1537_t) return std_logic_vector is
  variable rv : std_logic_vector(1536 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1537_t(x : std_logic_vector) return int1537_t is
  variable rv : int1537_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1538_t_to_slv(x : uint1538_t) return std_logic_vector is
  variable rv : std_logic_vector(1537 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1538_t(x : std_logic_vector) return uint1538_t is
  variable rv : uint1538_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1538_t_to_slv(x : int1538_t) return std_logic_vector is
  variable rv : std_logic_vector(1537 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1538_t(x : std_logic_vector) return int1538_t is
  variable rv : int1538_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1539_t_to_slv(x : uint1539_t) return std_logic_vector is
  variable rv : std_logic_vector(1538 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1539_t(x : std_logic_vector) return uint1539_t is
  variable rv : uint1539_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1539_t_to_slv(x : int1539_t) return std_logic_vector is
  variable rv : std_logic_vector(1538 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1539_t(x : std_logic_vector) return int1539_t is
  variable rv : int1539_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1540_t_to_slv(x : uint1540_t) return std_logic_vector is
  variable rv : std_logic_vector(1539 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1540_t(x : std_logic_vector) return uint1540_t is
  variable rv : uint1540_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1540_t_to_slv(x : int1540_t) return std_logic_vector is
  variable rv : std_logic_vector(1539 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1540_t(x : std_logic_vector) return int1540_t is
  variable rv : int1540_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1541_t_to_slv(x : uint1541_t) return std_logic_vector is
  variable rv : std_logic_vector(1540 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1541_t(x : std_logic_vector) return uint1541_t is
  variable rv : uint1541_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1541_t_to_slv(x : int1541_t) return std_logic_vector is
  variable rv : std_logic_vector(1540 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1541_t(x : std_logic_vector) return int1541_t is
  variable rv : int1541_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1542_t_to_slv(x : uint1542_t) return std_logic_vector is
  variable rv : std_logic_vector(1541 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1542_t(x : std_logic_vector) return uint1542_t is
  variable rv : uint1542_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1542_t_to_slv(x : int1542_t) return std_logic_vector is
  variable rv : std_logic_vector(1541 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1542_t(x : std_logic_vector) return int1542_t is
  variable rv : int1542_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1543_t_to_slv(x : uint1543_t) return std_logic_vector is
  variable rv : std_logic_vector(1542 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1543_t(x : std_logic_vector) return uint1543_t is
  variable rv : uint1543_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1543_t_to_slv(x : int1543_t) return std_logic_vector is
  variable rv : std_logic_vector(1542 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1543_t(x : std_logic_vector) return int1543_t is
  variable rv : int1543_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1544_t_to_slv(x : uint1544_t) return std_logic_vector is
  variable rv : std_logic_vector(1543 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1544_t(x : std_logic_vector) return uint1544_t is
  variable rv : uint1544_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1544_t_to_slv(x : int1544_t) return std_logic_vector is
  variable rv : std_logic_vector(1543 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1544_t(x : std_logic_vector) return int1544_t is
  variable rv : int1544_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1545_t_to_slv(x : uint1545_t) return std_logic_vector is
  variable rv : std_logic_vector(1544 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1545_t(x : std_logic_vector) return uint1545_t is
  variable rv : uint1545_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1545_t_to_slv(x : int1545_t) return std_logic_vector is
  variable rv : std_logic_vector(1544 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1545_t(x : std_logic_vector) return int1545_t is
  variable rv : int1545_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1546_t_to_slv(x : uint1546_t) return std_logic_vector is
  variable rv : std_logic_vector(1545 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1546_t(x : std_logic_vector) return uint1546_t is
  variable rv : uint1546_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1546_t_to_slv(x : int1546_t) return std_logic_vector is
  variable rv : std_logic_vector(1545 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1546_t(x : std_logic_vector) return int1546_t is
  variable rv : int1546_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1547_t_to_slv(x : uint1547_t) return std_logic_vector is
  variable rv : std_logic_vector(1546 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1547_t(x : std_logic_vector) return uint1547_t is
  variable rv : uint1547_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1547_t_to_slv(x : int1547_t) return std_logic_vector is
  variable rv : std_logic_vector(1546 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1547_t(x : std_logic_vector) return int1547_t is
  variable rv : int1547_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1548_t_to_slv(x : uint1548_t) return std_logic_vector is
  variable rv : std_logic_vector(1547 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1548_t(x : std_logic_vector) return uint1548_t is
  variable rv : uint1548_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1548_t_to_slv(x : int1548_t) return std_logic_vector is
  variable rv : std_logic_vector(1547 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1548_t(x : std_logic_vector) return int1548_t is
  variable rv : int1548_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1549_t_to_slv(x : uint1549_t) return std_logic_vector is
  variable rv : std_logic_vector(1548 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1549_t(x : std_logic_vector) return uint1549_t is
  variable rv : uint1549_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1549_t_to_slv(x : int1549_t) return std_logic_vector is
  variable rv : std_logic_vector(1548 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1549_t(x : std_logic_vector) return int1549_t is
  variable rv : int1549_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1550_t_to_slv(x : uint1550_t) return std_logic_vector is
  variable rv : std_logic_vector(1549 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1550_t(x : std_logic_vector) return uint1550_t is
  variable rv : uint1550_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1550_t_to_slv(x : int1550_t) return std_logic_vector is
  variable rv : std_logic_vector(1549 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1550_t(x : std_logic_vector) return int1550_t is
  variable rv : int1550_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1551_t_to_slv(x : uint1551_t) return std_logic_vector is
  variable rv : std_logic_vector(1550 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1551_t(x : std_logic_vector) return uint1551_t is
  variable rv : uint1551_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1551_t_to_slv(x : int1551_t) return std_logic_vector is
  variable rv : std_logic_vector(1550 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1551_t(x : std_logic_vector) return int1551_t is
  variable rv : int1551_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1552_t_to_slv(x : uint1552_t) return std_logic_vector is
  variable rv : std_logic_vector(1551 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1552_t(x : std_logic_vector) return uint1552_t is
  variable rv : uint1552_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1552_t_to_slv(x : int1552_t) return std_logic_vector is
  variable rv : std_logic_vector(1551 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1552_t(x : std_logic_vector) return int1552_t is
  variable rv : int1552_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1553_t_to_slv(x : uint1553_t) return std_logic_vector is
  variable rv : std_logic_vector(1552 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1553_t(x : std_logic_vector) return uint1553_t is
  variable rv : uint1553_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1553_t_to_slv(x : int1553_t) return std_logic_vector is
  variable rv : std_logic_vector(1552 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1553_t(x : std_logic_vector) return int1553_t is
  variable rv : int1553_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1554_t_to_slv(x : uint1554_t) return std_logic_vector is
  variable rv : std_logic_vector(1553 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1554_t(x : std_logic_vector) return uint1554_t is
  variable rv : uint1554_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1554_t_to_slv(x : int1554_t) return std_logic_vector is
  variable rv : std_logic_vector(1553 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1554_t(x : std_logic_vector) return int1554_t is
  variable rv : int1554_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1555_t_to_slv(x : uint1555_t) return std_logic_vector is
  variable rv : std_logic_vector(1554 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1555_t(x : std_logic_vector) return uint1555_t is
  variable rv : uint1555_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1555_t_to_slv(x : int1555_t) return std_logic_vector is
  variable rv : std_logic_vector(1554 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1555_t(x : std_logic_vector) return int1555_t is
  variable rv : int1555_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1556_t_to_slv(x : uint1556_t) return std_logic_vector is
  variable rv : std_logic_vector(1555 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1556_t(x : std_logic_vector) return uint1556_t is
  variable rv : uint1556_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1556_t_to_slv(x : int1556_t) return std_logic_vector is
  variable rv : std_logic_vector(1555 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1556_t(x : std_logic_vector) return int1556_t is
  variable rv : int1556_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1557_t_to_slv(x : uint1557_t) return std_logic_vector is
  variable rv : std_logic_vector(1556 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1557_t(x : std_logic_vector) return uint1557_t is
  variable rv : uint1557_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1557_t_to_slv(x : int1557_t) return std_logic_vector is
  variable rv : std_logic_vector(1556 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1557_t(x : std_logic_vector) return int1557_t is
  variable rv : int1557_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1558_t_to_slv(x : uint1558_t) return std_logic_vector is
  variable rv : std_logic_vector(1557 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1558_t(x : std_logic_vector) return uint1558_t is
  variable rv : uint1558_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1558_t_to_slv(x : int1558_t) return std_logic_vector is
  variable rv : std_logic_vector(1557 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1558_t(x : std_logic_vector) return int1558_t is
  variable rv : int1558_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1559_t_to_slv(x : uint1559_t) return std_logic_vector is
  variable rv : std_logic_vector(1558 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1559_t(x : std_logic_vector) return uint1559_t is
  variable rv : uint1559_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1559_t_to_slv(x : int1559_t) return std_logic_vector is
  variable rv : std_logic_vector(1558 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1559_t(x : std_logic_vector) return int1559_t is
  variable rv : int1559_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1560_t_to_slv(x : uint1560_t) return std_logic_vector is
  variable rv : std_logic_vector(1559 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1560_t(x : std_logic_vector) return uint1560_t is
  variable rv : uint1560_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1560_t_to_slv(x : int1560_t) return std_logic_vector is
  variable rv : std_logic_vector(1559 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1560_t(x : std_logic_vector) return int1560_t is
  variable rv : int1560_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1561_t_to_slv(x : uint1561_t) return std_logic_vector is
  variable rv : std_logic_vector(1560 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1561_t(x : std_logic_vector) return uint1561_t is
  variable rv : uint1561_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1561_t_to_slv(x : int1561_t) return std_logic_vector is
  variable rv : std_logic_vector(1560 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1561_t(x : std_logic_vector) return int1561_t is
  variable rv : int1561_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1562_t_to_slv(x : uint1562_t) return std_logic_vector is
  variable rv : std_logic_vector(1561 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1562_t(x : std_logic_vector) return uint1562_t is
  variable rv : uint1562_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1562_t_to_slv(x : int1562_t) return std_logic_vector is
  variable rv : std_logic_vector(1561 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1562_t(x : std_logic_vector) return int1562_t is
  variable rv : int1562_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1563_t_to_slv(x : uint1563_t) return std_logic_vector is
  variable rv : std_logic_vector(1562 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1563_t(x : std_logic_vector) return uint1563_t is
  variable rv : uint1563_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1563_t_to_slv(x : int1563_t) return std_logic_vector is
  variable rv : std_logic_vector(1562 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1563_t(x : std_logic_vector) return int1563_t is
  variable rv : int1563_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1564_t_to_slv(x : uint1564_t) return std_logic_vector is
  variable rv : std_logic_vector(1563 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1564_t(x : std_logic_vector) return uint1564_t is
  variable rv : uint1564_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1564_t_to_slv(x : int1564_t) return std_logic_vector is
  variable rv : std_logic_vector(1563 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1564_t(x : std_logic_vector) return int1564_t is
  variable rv : int1564_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1565_t_to_slv(x : uint1565_t) return std_logic_vector is
  variable rv : std_logic_vector(1564 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1565_t(x : std_logic_vector) return uint1565_t is
  variable rv : uint1565_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1565_t_to_slv(x : int1565_t) return std_logic_vector is
  variable rv : std_logic_vector(1564 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1565_t(x : std_logic_vector) return int1565_t is
  variable rv : int1565_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1566_t_to_slv(x : uint1566_t) return std_logic_vector is
  variable rv : std_logic_vector(1565 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1566_t(x : std_logic_vector) return uint1566_t is
  variable rv : uint1566_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1566_t_to_slv(x : int1566_t) return std_logic_vector is
  variable rv : std_logic_vector(1565 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1566_t(x : std_logic_vector) return int1566_t is
  variable rv : int1566_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1567_t_to_slv(x : uint1567_t) return std_logic_vector is
  variable rv : std_logic_vector(1566 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1567_t(x : std_logic_vector) return uint1567_t is
  variable rv : uint1567_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1567_t_to_slv(x : int1567_t) return std_logic_vector is
  variable rv : std_logic_vector(1566 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1567_t(x : std_logic_vector) return int1567_t is
  variable rv : int1567_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1568_t_to_slv(x : uint1568_t) return std_logic_vector is
  variable rv : std_logic_vector(1567 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1568_t(x : std_logic_vector) return uint1568_t is
  variable rv : uint1568_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1568_t_to_slv(x : int1568_t) return std_logic_vector is
  variable rv : std_logic_vector(1567 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1568_t(x : std_logic_vector) return int1568_t is
  variable rv : int1568_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1569_t_to_slv(x : uint1569_t) return std_logic_vector is
  variable rv : std_logic_vector(1568 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1569_t(x : std_logic_vector) return uint1569_t is
  variable rv : uint1569_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1569_t_to_slv(x : int1569_t) return std_logic_vector is
  variable rv : std_logic_vector(1568 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1569_t(x : std_logic_vector) return int1569_t is
  variable rv : int1569_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1570_t_to_slv(x : uint1570_t) return std_logic_vector is
  variable rv : std_logic_vector(1569 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1570_t(x : std_logic_vector) return uint1570_t is
  variable rv : uint1570_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1570_t_to_slv(x : int1570_t) return std_logic_vector is
  variable rv : std_logic_vector(1569 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1570_t(x : std_logic_vector) return int1570_t is
  variable rv : int1570_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1571_t_to_slv(x : uint1571_t) return std_logic_vector is
  variable rv : std_logic_vector(1570 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1571_t(x : std_logic_vector) return uint1571_t is
  variable rv : uint1571_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1571_t_to_slv(x : int1571_t) return std_logic_vector is
  variable rv : std_logic_vector(1570 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1571_t(x : std_logic_vector) return int1571_t is
  variable rv : int1571_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1572_t_to_slv(x : uint1572_t) return std_logic_vector is
  variable rv : std_logic_vector(1571 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1572_t(x : std_logic_vector) return uint1572_t is
  variable rv : uint1572_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1572_t_to_slv(x : int1572_t) return std_logic_vector is
  variable rv : std_logic_vector(1571 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1572_t(x : std_logic_vector) return int1572_t is
  variable rv : int1572_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1573_t_to_slv(x : uint1573_t) return std_logic_vector is
  variable rv : std_logic_vector(1572 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1573_t(x : std_logic_vector) return uint1573_t is
  variable rv : uint1573_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1573_t_to_slv(x : int1573_t) return std_logic_vector is
  variable rv : std_logic_vector(1572 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1573_t(x : std_logic_vector) return int1573_t is
  variable rv : int1573_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1574_t_to_slv(x : uint1574_t) return std_logic_vector is
  variable rv : std_logic_vector(1573 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1574_t(x : std_logic_vector) return uint1574_t is
  variable rv : uint1574_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1574_t_to_slv(x : int1574_t) return std_logic_vector is
  variable rv : std_logic_vector(1573 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1574_t(x : std_logic_vector) return int1574_t is
  variable rv : int1574_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1575_t_to_slv(x : uint1575_t) return std_logic_vector is
  variable rv : std_logic_vector(1574 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1575_t(x : std_logic_vector) return uint1575_t is
  variable rv : uint1575_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1575_t_to_slv(x : int1575_t) return std_logic_vector is
  variable rv : std_logic_vector(1574 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1575_t(x : std_logic_vector) return int1575_t is
  variable rv : int1575_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1576_t_to_slv(x : uint1576_t) return std_logic_vector is
  variable rv : std_logic_vector(1575 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1576_t(x : std_logic_vector) return uint1576_t is
  variable rv : uint1576_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1576_t_to_slv(x : int1576_t) return std_logic_vector is
  variable rv : std_logic_vector(1575 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1576_t(x : std_logic_vector) return int1576_t is
  variable rv : int1576_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1577_t_to_slv(x : uint1577_t) return std_logic_vector is
  variable rv : std_logic_vector(1576 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1577_t(x : std_logic_vector) return uint1577_t is
  variable rv : uint1577_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1577_t_to_slv(x : int1577_t) return std_logic_vector is
  variable rv : std_logic_vector(1576 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1577_t(x : std_logic_vector) return int1577_t is
  variable rv : int1577_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1578_t_to_slv(x : uint1578_t) return std_logic_vector is
  variable rv : std_logic_vector(1577 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1578_t(x : std_logic_vector) return uint1578_t is
  variable rv : uint1578_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1578_t_to_slv(x : int1578_t) return std_logic_vector is
  variable rv : std_logic_vector(1577 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1578_t(x : std_logic_vector) return int1578_t is
  variable rv : int1578_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1579_t_to_slv(x : uint1579_t) return std_logic_vector is
  variable rv : std_logic_vector(1578 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1579_t(x : std_logic_vector) return uint1579_t is
  variable rv : uint1579_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1579_t_to_slv(x : int1579_t) return std_logic_vector is
  variable rv : std_logic_vector(1578 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1579_t(x : std_logic_vector) return int1579_t is
  variable rv : int1579_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1580_t_to_slv(x : uint1580_t) return std_logic_vector is
  variable rv : std_logic_vector(1579 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1580_t(x : std_logic_vector) return uint1580_t is
  variable rv : uint1580_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1580_t_to_slv(x : int1580_t) return std_logic_vector is
  variable rv : std_logic_vector(1579 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1580_t(x : std_logic_vector) return int1580_t is
  variable rv : int1580_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1581_t_to_slv(x : uint1581_t) return std_logic_vector is
  variable rv : std_logic_vector(1580 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1581_t(x : std_logic_vector) return uint1581_t is
  variable rv : uint1581_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1581_t_to_slv(x : int1581_t) return std_logic_vector is
  variable rv : std_logic_vector(1580 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1581_t(x : std_logic_vector) return int1581_t is
  variable rv : int1581_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1582_t_to_slv(x : uint1582_t) return std_logic_vector is
  variable rv : std_logic_vector(1581 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1582_t(x : std_logic_vector) return uint1582_t is
  variable rv : uint1582_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1582_t_to_slv(x : int1582_t) return std_logic_vector is
  variable rv : std_logic_vector(1581 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1582_t(x : std_logic_vector) return int1582_t is
  variable rv : int1582_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1583_t_to_slv(x : uint1583_t) return std_logic_vector is
  variable rv : std_logic_vector(1582 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1583_t(x : std_logic_vector) return uint1583_t is
  variable rv : uint1583_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1583_t_to_slv(x : int1583_t) return std_logic_vector is
  variable rv : std_logic_vector(1582 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1583_t(x : std_logic_vector) return int1583_t is
  variable rv : int1583_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1584_t_to_slv(x : uint1584_t) return std_logic_vector is
  variable rv : std_logic_vector(1583 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1584_t(x : std_logic_vector) return uint1584_t is
  variable rv : uint1584_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1584_t_to_slv(x : int1584_t) return std_logic_vector is
  variable rv : std_logic_vector(1583 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1584_t(x : std_logic_vector) return int1584_t is
  variable rv : int1584_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1585_t_to_slv(x : uint1585_t) return std_logic_vector is
  variable rv : std_logic_vector(1584 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1585_t(x : std_logic_vector) return uint1585_t is
  variable rv : uint1585_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1585_t_to_slv(x : int1585_t) return std_logic_vector is
  variable rv : std_logic_vector(1584 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1585_t(x : std_logic_vector) return int1585_t is
  variable rv : int1585_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1586_t_to_slv(x : uint1586_t) return std_logic_vector is
  variable rv : std_logic_vector(1585 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1586_t(x : std_logic_vector) return uint1586_t is
  variable rv : uint1586_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1586_t_to_slv(x : int1586_t) return std_logic_vector is
  variable rv : std_logic_vector(1585 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1586_t(x : std_logic_vector) return int1586_t is
  variable rv : int1586_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1587_t_to_slv(x : uint1587_t) return std_logic_vector is
  variable rv : std_logic_vector(1586 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1587_t(x : std_logic_vector) return uint1587_t is
  variable rv : uint1587_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1587_t_to_slv(x : int1587_t) return std_logic_vector is
  variable rv : std_logic_vector(1586 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1587_t(x : std_logic_vector) return int1587_t is
  variable rv : int1587_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1588_t_to_slv(x : uint1588_t) return std_logic_vector is
  variable rv : std_logic_vector(1587 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1588_t(x : std_logic_vector) return uint1588_t is
  variable rv : uint1588_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1588_t_to_slv(x : int1588_t) return std_logic_vector is
  variable rv : std_logic_vector(1587 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1588_t(x : std_logic_vector) return int1588_t is
  variable rv : int1588_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1589_t_to_slv(x : uint1589_t) return std_logic_vector is
  variable rv : std_logic_vector(1588 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1589_t(x : std_logic_vector) return uint1589_t is
  variable rv : uint1589_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1589_t_to_slv(x : int1589_t) return std_logic_vector is
  variable rv : std_logic_vector(1588 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1589_t(x : std_logic_vector) return int1589_t is
  variable rv : int1589_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1590_t_to_slv(x : uint1590_t) return std_logic_vector is
  variable rv : std_logic_vector(1589 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1590_t(x : std_logic_vector) return uint1590_t is
  variable rv : uint1590_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1590_t_to_slv(x : int1590_t) return std_logic_vector is
  variable rv : std_logic_vector(1589 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1590_t(x : std_logic_vector) return int1590_t is
  variable rv : int1590_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1591_t_to_slv(x : uint1591_t) return std_logic_vector is
  variable rv : std_logic_vector(1590 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1591_t(x : std_logic_vector) return uint1591_t is
  variable rv : uint1591_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1591_t_to_slv(x : int1591_t) return std_logic_vector is
  variable rv : std_logic_vector(1590 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1591_t(x : std_logic_vector) return int1591_t is
  variable rv : int1591_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1592_t_to_slv(x : uint1592_t) return std_logic_vector is
  variable rv : std_logic_vector(1591 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1592_t(x : std_logic_vector) return uint1592_t is
  variable rv : uint1592_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1592_t_to_slv(x : int1592_t) return std_logic_vector is
  variable rv : std_logic_vector(1591 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1592_t(x : std_logic_vector) return int1592_t is
  variable rv : int1592_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1593_t_to_slv(x : uint1593_t) return std_logic_vector is
  variable rv : std_logic_vector(1592 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1593_t(x : std_logic_vector) return uint1593_t is
  variable rv : uint1593_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1593_t_to_slv(x : int1593_t) return std_logic_vector is
  variable rv : std_logic_vector(1592 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1593_t(x : std_logic_vector) return int1593_t is
  variable rv : int1593_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1594_t_to_slv(x : uint1594_t) return std_logic_vector is
  variable rv : std_logic_vector(1593 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1594_t(x : std_logic_vector) return uint1594_t is
  variable rv : uint1594_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1594_t_to_slv(x : int1594_t) return std_logic_vector is
  variable rv : std_logic_vector(1593 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1594_t(x : std_logic_vector) return int1594_t is
  variable rv : int1594_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1595_t_to_slv(x : uint1595_t) return std_logic_vector is
  variable rv : std_logic_vector(1594 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1595_t(x : std_logic_vector) return uint1595_t is
  variable rv : uint1595_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1595_t_to_slv(x : int1595_t) return std_logic_vector is
  variable rv : std_logic_vector(1594 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1595_t(x : std_logic_vector) return int1595_t is
  variable rv : int1595_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1596_t_to_slv(x : uint1596_t) return std_logic_vector is
  variable rv : std_logic_vector(1595 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1596_t(x : std_logic_vector) return uint1596_t is
  variable rv : uint1596_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1596_t_to_slv(x : int1596_t) return std_logic_vector is
  variable rv : std_logic_vector(1595 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1596_t(x : std_logic_vector) return int1596_t is
  variable rv : int1596_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1597_t_to_slv(x : uint1597_t) return std_logic_vector is
  variable rv : std_logic_vector(1596 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1597_t(x : std_logic_vector) return uint1597_t is
  variable rv : uint1597_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1597_t_to_slv(x : int1597_t) return std_logic_vector is
  variable rv : std_logic_vector(1596 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1597_t(x : std_logic_vector) return int1597_t is
  variable rv : int1597_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1598_t_to_slv(x : uint1598_t) return std_logic_vector is
  variable rv : std_logic_vector(1597 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1598_t(x : std_logic_vector) return uint1598_t is
  variable rv : uint1598_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1598_t_to_slv(x : int1598_t) return std_logic_vector is
  variable rv : std_logic_vector(1597 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1598_t(x : std_logic_vector) return int1598_t is
  variable rv : int1598_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1599_t_to_slv(x : uint1599_t) return std_logic_vector is
  variable rv : std_logic_vector(1598 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1599_t(x : std_logic_vector) return uint1599_t is
  variable rv : uint1599_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1599_t_to_slv(x : int1599_t) return std_logic_vector is
  variable rv : std_logic_vector(1598 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1599_t(x : std_logic_vector) return int1599_t is
  variable rv : int1599_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1600_t_to_slv(x : uint1600_t) return std_logic_vector is
  variable rv : std_logic_vector(1599 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1600_t(x : std_logic_vector) return uint1600_t is
  variable rv : uint1600_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1600_t_to_slv(x : int1600_t) return std_logic_vector is
  variable rv : std_logic_vector(1599 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1600_t(x : std_logic_vector) return int1600_t is
  variable rv : int1600_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1601_t_to_slv(x : uint1601_t) return std_logic_vector is
  variable rv : std_logic_vector(1600 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1601_t(x : std_logic_vector) return uint1601_t is
  variable rv : uint1601_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1601_t_to_slv(x : int1601_t) return std_logic_vector is
  variable rv : std_logic_vector(1600 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1601_t(x : std_logic_vector) return int1601_t is
  variable rv : int1601_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1602_t_to_slv(x : uint1602_t) return std_logic_vector is
  variable rv : std_logic_vector(1601 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1602_t(x : std_logic_vector) return uint1602_t is
  variable rv : uint1602_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1602_t_to_slv(x : int1602_t) return std_logic_vector is
  variable rv : std_logic_vector(1601 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1602_t(x : std_logic_vector) return int1602_t is
  variable rv : int1602_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1603_t_to_slv(x : uint1603_t) return std_logic_vector is
  variable rv : std_logic_vector(1602 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1603_t(x : std_logic_vector) return uint1603_t is
  variable rv : uint1603_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1603_t_to_slv(x : int1603_t) return std_logic_vector is
  variable rv : std_logic_vector(1602 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1603_t(x : std_logic_vector) return int1603_t is
  variable rv : int1603_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1604_t_to_slv(x : uint1604_t) return std_logic_vector is
  variable rv : std_logic_vector(1603 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1604_t(x : std_logic_vector) return uint1604_t is
  variable rv : uint1604_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1604_t_to_slv(x : int1604_t) return std_logic_vector is
  variable rv : std_logic_vector(1603 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1604_t(x : std_logic_vector) return int1604_t is
  variable rv : int1604_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1605_t_to_slv(x : uint1605_t) return std_logic_vector is
  variable rv : std_logic_vector(1604 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1605_t(x : std_logic_vector) return uint1605_t is
  variable rv : uint1605_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1605_t_to_slv(x : int1605_t) return std_logic_vector is
  variable rv : std_logic_vector(1604 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1605_t(x : std_logic_vector) return int1605_t is
  variable rv : int1605_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1606_t_to_slv(x : uint1606_t) return std_logic_vector is
  variable rv : std_logic_vector(1605 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1606_t(x : std_logic_vector) return uint1606_t is
  variable rv : uint1606_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1606_t_to_slv(x : int1606_t) return std_logic_vector is
  variable rv : std_logic_vector(1605 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1606_t(x : std_logic_vector) return int1606_t is
  variable rv : int1606_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1607_t_to_slv(x : uint1607_t) return std_logic_vector is
  variable rv : std_logic_vector(1606 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1607_t(x : std_logic_vector) return uint1607_t is
  variable rv : uint1607_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1607_t_to_slv(x : int1607_t) return std_logic_vector is
  variable rv : std_logic_vector(1606 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1607_t(x : std_logic_vector) return int1607_t is
  variable rv : int1607_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1608_t_to_slv(x : uint1608_t) return std_logic_vector is
  variable rv : std_logic_vector(1607 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1608_t(x : std_logic_vector) return uint1608_t is
  variable rv : uint1608_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1608_t_to_slv(x : int1608_t) return std_logic_vector is
  variable rv : std_logic_vector(1607 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1608_t(x : std_logic_vector) return int1608_t is
  variable rv : int1608_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1609_t_to_slv(x : uint1609_t) return std_logic_vector is
  variable rv : std_logic_vector(1608 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1609_t(x : std_logic_vector) return uint1609_t is
  variable rv : uint1609_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1609_t_to_slv(x : int1609_t) return std_logic_vector is
  variable rv : std_logic_vector(1608 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1609_t(x : std_logic_vector) return int1609_t is
  variable rv : int1609_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1610_t_to_slv(x : uint1610_t) return std_logic_vector is
  variable rv : std_logic_vector(1609 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1610_t(x : std_logic_vector) return uint1610_t is
  variable rv : uint1610_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1610_t_to_slv(x : int1610_t) return std_logic_vector is
  variable rv : std_logic_vector(1609 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1610_t(x : std_logic_vector) return int1610_t is
  variable rv : int1610_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1611_t_to_slv(x : uint1611_t) return std_logic_vector is
  variable rv : std_logic_vector(1610 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1611_t(x : std_logic_vector) return uint1611_t is
  variable rv : uint1611_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1611_t_to_slv(x : int1611_t) return std_logic_vector is
  variable rv : std_logic_vector(1610 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1611_t(x : std_logic_vector) return int1611_t is
  variable rv : int1611_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1612_t_to_slv(x : uint1612_t) return std_logic_vector is
  variable rv : std_logic_vector(1611 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1612_t(x : std_logic_vector) return uint1612_t is
  variable rv : uint1612_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1612_t_to_slv(x : int1612_t) return std_logic_vector is
  variable rv : std_logic_vector(1611 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1612_t(x : std_logic_vector) return int1612_t is
  variable rv : int1612_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1613_t_to_slv(x : uint1613_t) return std_logic_vector is
  variable rv : std_logic_vector(1612 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1613_t(x : std_logic_vector) return uint1613_t is
  variable rv : uint1613_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1613_t_to_slv(x : int1613_t) return std_logic_vector is
  variable rv : std_logic_vector(1612 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1613_t(x : std_logic_vector) return int1613_t is
  variable rv : int1613_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1614_t_to_slv(x : uint1614_t) return std_logic_vector is
  variable rv : std_logic_vector(1613 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1614_t(x : std_logic_vector) return uint1614_t is
  variable rv : uint1614_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1614_t_to_slv(x : int1614_t) return std_logic_vector is
  variable rv : std_logic_vector(1613 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1614_t(x : std_logic_vector) return int1614_t is
  variable rv : int1614_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1615_t_to_slv(x : uint1615_t) return std_logic_vector is
  variable rv : std_logic_vector(1614 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1615_t(x : std_logic_vector) return uint1615_t is
  variable rv : uint1615_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1615_t_to_slv(x : int1615_t) return std_logic_vector is
  variable rv : std_logic_vector(1614 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1615_t(x : std_logic_vector) return int1615_t is
  variable rv : int1615_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1616_t_to_slv(x : uint1616_t) return std_logic_vector is
  variable rv : std_logic_vector(1615 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1616_t(x : std_logic_vector) return uint1616_t is
  variable rv : uint1616_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1616_t_to_slv(x : int1616_t) return std_logic_vector is
  variable rv : std_logic_vector(1615 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1616_t(x : std_logic_vector) return int1616_t is
  variable rv : int1616_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1617_t_to_slv(x : uint1617_t) return std_logic_vector is
  variable rv : std_logic_vector(1616 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1617_t(x : std_logic_vector) return uint1617_t is
  variable rv : uint1617_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1617_t_to_slv(x : int1617_t) return std_logic_vector is
  variable rv : std_logic_vector(1616 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1617_t(x : std_logic_vector) return int1617_t is
  variable rv : int1617_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1618_t_to_slv(x : uint1618_t) return std_logic_vector is
  variable rv : std_logic_vector(1617 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1618_t(x : std_logic_vector) return uint1618_t is
  variable rv : uint1618_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1618_t_to_slv(x : int1618_t) return std_logic_vector is
  variable rv : std_logic_vector(1617 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1618_t(x : std_logic_vector) return int1618_t is
  variable rv : int1618_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1619_t_to_slv(x : uint1619_t) return std_logic_vector is
  variable rv : std_logic_vector(1618 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1619_t(x : std_logic_vector) return uint1619_t is
  variable rv : uint1619_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1619_t_to_slv(x : int1619_t) return std_logic_vector is
  variable rv : std_logic_vector(1618 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1619_t(x : std_logic_vector) return int1619_t is
  variable rv : int1619_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1620_t_to_slv(x : uint1620_t) return std_logic_vector is
  variable rv : std_logic_vector(1619 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1620_t(x : std_logic_vector) return uint1620_t is
  variable rv : uint1620_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1620_t_to_slv(x : int1620_t) return std_logic_vector is
  variable rv : std_logic_vector(1619 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1620_t(x : std_logic_vector) return int1620_t is
  variable rv : int1620_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1621_t_to_slv(x : uint1621_t) return std_logic_vector is
  variable rv : std_logic_vector(1620 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1621_t(x : std_logic_vector) return uint1621_t is
  variable rv : uint1621_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1621_t_to_slv(x : int1621_t) return std_logic_vector is
  variable rv : std_logic_vector(1620 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1621_t(x : std_logic_vector) return int1621_t is
  variable rv : int1621_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1622_t_to_slv(x : uint1622_t) return std_logic_vector is
  variable rv : std_logic_vector(1621 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1622_t(x : std_logic_vector) return uint1622_t is
  variable rv : uint1622_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1622_t_to_slv(x : int1622_t) return std_logic_vector is
  variable rv : std_logic_vector(1621 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1622_t(x : std_logic_vector) return int1622_t is
  variable rv : int1622_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1623_t_to_slv(x : uint1623_t) return std_logic_vector is
  variable rv : std_logic_vector(1622 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1623_t(x : std_logic_vector) return uint1623_t is
  variable rv : uint1623_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1623_t_to_slv(x : int1623_t) return std_logic_vector is
  variable rv : std_logic_vector(1622 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1623_t(x : std_logic_vector) return int1623_t is
  variable rv : int1623_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1624_t_to_slv(x : uint1624_t) return std_logic_vector is
  variable rv : std_logic_vector(1623 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1624_t(x : std_logic_vector) return uint1624_t is
  variable rv : uint1624_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1624_t_to_slv(x : int1624_t) return std_logic_vector is
  variable rv : std_logic_vector(1623 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1624_t(x : std_logic_vector) return int1624_t is
  variable rv : int1624_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1625_t_to_slv(x : uint1625_t) return std_logic_vector is
  variable rv : std_logic_vector(1624 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1625_t(x : std_logic_vector) return uint1625_t is
  variable rv : uint1625_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1625_t_to_slv(x : int1625_t) return std_logic_vector is
  variable rv : std_logic_vector(1624 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1625_t(x : std_logic_vector) return int1625_t is
  variable rv : int1625_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1626_t_to_slv(x : uint1626_t) return std_logic_vector is
  variable rv : std_logic_vector(1625 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1626_t(x : std_logic_vector) return uint1626_t is
  variable rv : uint1626_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1626_t_to_slv(x : int1626_t) return std_logic_vector is
  variable rv : std_logic_vector(1625 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1626_t(x : std_logic_vector) return int1626_t is
  variable rv : int1626_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1627_t_to_slv(x : uint1627_t) return std_logic_vector is
  variable rv : std_logic_vector(1626 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1627_t(x : std_logic_vector) return uint1627_t is
  variable rv : uint1627_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1627_t_to_slv(x : int1627_t) return std_logic_vector is
  variable rv : std_logic_vector(1626 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1627_t(x : std_logic_vector) return int1627_t is
  variable rv : int1627_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1628_t_to_slv(x : uint1628_t) return std_logic_vector is
  variable rv : std_logic_vector(1627 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1628_t(x : std_logic_vector) return uint1628_t is
  variable rv : uint1628_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1628_t_to_slv(x : int1628_t) return std_logic_vector is
  variable rv : std_logic_vector(1627 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1628_t(x : std_logic_vector) return int1628_t is
  variable rv : int1628_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1629_t_to_slv(x : uint1629_t) return std_logic_vector is
  variable rv : std_logic_vector(1628 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1629_t(x : std_logic_vector) return uint1629_t is
  variable rv : uint1629_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1629_t_to_slv(x : int1629_t) return std_logic_vector is
  variable rv : std_logic_vector(1628 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1629_t(x : std_logic_vector) return int1629_t is
  variable rv : int1629_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1630_t_to_slv(x : uint1630_t) return std_logic_vector is
  variable rv : std_logic_vector(1629 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1630_t(x : std_logic_vector) return uint1630_t is
  variable rv : uint1630_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1630_t_to_slv(x : int1630_t) return std_logic_vector is
  variable rv : std_logic_vector(1629 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1630_t(x : std_logic_vector) return int1630_t is
  variable rv : int1630_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1631_t_to_slv(x : uint1631_t) return std_logic_vector is
  variable rv : std_logic_vector(1630 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1631_t(x : std_logic_vector) return uint1631_t is
  variable rv : uint1631_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1631_t_to_slv(x : int1631_t) return std_logic_vector is
  variable rv : std_logic_vector(1630 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1631_t(x : std_logic_vector) return int1631_t is
  variable rv : int1631_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1632_t_to_slv(x : uint1632_t) return std_logic_vector is
  variable rv : std_logic_vector(1631 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1632_t(x : std_logic_vector) return uint1632_t is
  variable rv : uint1632_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1632_t_to_slv(x : int1632_t) return std_logic_vector is
  variable rv : std_logic_vector(1631 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1632_t(x : std_logic_vector) return int1632_t is
  variable rv : int1632_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1633_t_to_slv(x : uint1633_t) return std_logic_vector is
  variable rv : std_logic_vector(1632 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1633_t(x : std_logic_vector) return uint1633_t is
  variable rv : uint1633_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1633_t_to_slv(x : int1633_t) return std_logic_vector is
  variable rv : std_logic_vector(1632 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1633_t(x : std_logic_vector) return int1633_t is
  variable rv : int1633_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1634_t_to_slv(x : uint1634_t) return std_logic_vector is
  variable rv : std_logic_vector(1633 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1634_t(x : std_logic_vector) return uint1634_t is
  variable rv : uint1634_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1634_t_to_slv(x : int1634_t) return std_logic_vector is
  variable rv : std_logic_vector(1633 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1634_t(x : std_logic_vector) return int1634_t is
  variable rv : int1634_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1635_t_to_slv(x : uint1635_t) return std_logic_vector is
  variable rv : std_logic_vector(1634 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1635_t(x : std_logic_vector) return uint1635_t is
  variable rv : uint1635_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1635_t_to_slv(x : int1635_t) return std_logic_vector is
  variable rv : std_logic_vector(1634 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1635_t(x : std_logic_vector) return int1635_t is
  variable rv : int1635_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1636_t_to_slv(x : uint1636_t) return std_logic_vector is
  variable rv : std_logic_vector(1635 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1636_t(x : std_logic_vector) return uint1636_t is
  variable rv : uint1636_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1636_t_to_slv(x : int1636_t) return std_logic_vector is
  variable rv : std_logic_vector(1635 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1636_t(x : std_logic_vector) return int1636_t is
  variable rv : int1636_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1637_t_to_slv(x : uint1637_t) return std_logic_vector is
  variable rv : std_logic_vector(1636 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1637_t(x : std_logic_vector) return uint1637_t is
  variable rv : uint1637_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1637_t_to_slv(x : int1637_t) return std_logic_vector is
  variable rv : std_logic_vector(1636 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1637_t(x : std_logic_vector) return int1637_t is
  variable rv : int1637_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1638_t_to_slv(x : uint1638_t) return std_logic_vector is
  variable rv : std_logic_vector(1637 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1638_t(x : std_logic_vector) return uint1638_t is
  variable rv : uint1638_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1638_t_to_slv(x : int1638_t) return std_logic_vector is
  variable rv : std_logic_vector(1637 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1638_t(x : std_logic_vector) return int1638_t is
  variable rv : int1638_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1639_t_to_slv(x : uint1639_t) return std_logic_vector is
  variable rv : std_logic_vector(1638 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1639_t(x : std_logic_vector) return uint1639_t is
  variable rv : uint1639_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1639_t_to_slv(x : int1639_t) return std_logic_vector is
  variable rv : std_logic_vector(1638 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1639_t(x : std_logic_vector) return int1639_t is
  variable rv : int1639_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1640_t_to_slv(x : uint1640_t) return std_logic_vector is
  variable rv : std_logic_vector(1639 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1640_t(x : std_logic_vector) return uint1640_t is
  variable rv : uint1640_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1640_t_to_slv(x : int1640_t) return std_logic_vector is
  variable rv : std_logic_vector(1639 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1640_t(x : std_logic_vector) return int1640_t is
  variable rv : int1640_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1641_t_to_slv(x : uint1641_t) return std_logic_vector is
  variable rv : std_logic_vector(1640 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1641_t(x : std_logic_vector) return uint1641_t is
  variable rv : uint1641_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1641_t_to_slv(x : int1641_t) return std_logic_vector is
  variable rv : std_logic_vector(1640 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1641_t(x : std_logic_vector) return int1641_t is
  variable rv : int1641_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1642_t_to_slv(x : uint1642_t) return std_logic_vector is
  variable rv : std_logic_vector(1641 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1642_t(x : std_logic_vector) return uint1642_t is
  variable rv : uint1642_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1642_t_to_slv(x : int1642_t) return std_logic_vector is
  variable rv : std_logic_vector(1641 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1642_t(x : std_logic_vector) return int1642_t is
  variable rv : int1642_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1643_t_to_slv(x : uint1643_t) return std_logic_vector is
  variable rv : std_logic_vector(1642 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1643_t(x : std_logic_vector) return uint1643_t is
  variable rv : uint1643_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1643_t_to_slv(x : int1643_t) return std_logic_vector is
  variable rv : std_logic_vector(1642 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1643_t(x : std_logic_vector) return int1643_t is
  variable rv : int1643_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1644_t_to_slv(x : uint1644_t) return std_logic_vector is
  variable rv : std_logic_vector(1643 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1644_t(x : std_logic_vector) return uint1644_t is
  variable rv : uint1644_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1644_t_to_slv(x : int1644_t) return std_logic_vector is
  variable rv : std_logic_vector(1643 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1644_t(x : std_logic_vector) return int1644_t is
  variable rv : int1644_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1645_t_to_slv(x : uint1645_t) return std_logic_vector is
  variable rv : std_logic_vector(1644 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1645_t(x : std_logic_vector) return uint1645_t is
  variable rv : uint1645_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1645_t_to_slv(x : int1645_t) return std_logic_vector is
  variable rv : std_logic_vector(1644 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1645_t(x : std_logic_vector) return int1645_t is
  variable rv : int1645_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1646_t_to_slv(x : uint1646_t) return std_logic_vector is
  variable rv : std_logic_vector(1645 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1646_t(x : std_logic_vector) return uint1646_t is
  variable rv : uint1646_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1646_t_to_slv(x : int1646_t) return std_logic_vector is
  variable rv : std_logic_vector(1645 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1646_t(x : std_logic_vector) return int1646_t is
  variable rv : int1646_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1647_t_to_slv(x : uint1647_t) return std_logic_vector is
  variable rv : std_logic_vector(1646 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1647_t(x : std_logic_vector) return uint1647_t is
  variable rv : uint1647_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1647_t_to_slv(x : int1647_t) return std_logic_vector is
  variable rv : std_logic_vector(1646 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1647_t(x : std_logic_vector) return int1647_t is
  variable rv : int1647_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1648_t_to_slv(x : uint1648_t) return std_logic_vector is
  variable rv : std_logic_vector(1647 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1648_t(x : std_logic_vector) return uint1648_t is
  variable rv : uint1648_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1648_t_to_slv(x : int1648_t) return std_logic_vector is
  variable rv : std_logic_vector(1647 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1648_t(x : std_logic_vector) return int1648_t is
  variable rv : int1648_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1649_t_to_slv(x : uint1649_t) return std_logic_vector is
  variable rv : std_logic_vector(1648 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1649_t(x : std_logic_vector) return uint1649_t is
  variable rv : uint1649_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1649_t_to_slv(x : int1649_t) return std_logic_vector is
  variable rv : std_logic_vector(1648 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1649_t(x : std_logic_vector) return int1649_t is
  variable rv : int1649_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1650_t_to_slv(x : uint1650_t) return std_logic_vector is
  variable rv : std_logic_vector(1649 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1650_t(x : std_logic_vector) return uint1650_t is
  variable rv : uint1650_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1650_t_to_slv(x : int1650_t) return std_logic_vector is
  variable rv : std_logic_vector(1649 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1650_t(x : std_logic_vector) return int1650_t is
  variable rv : int1650_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1651_t_to_slv(x : uint1651_t) return std_logic_vector is
  variable rv : std_logic_vector(1650 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1651_t(x : std_logic_vector) return uint1651_t is
  variable rv : uint1651_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1651_t_to_slv(x : int1651_t) return std_logic_vector is
  variable rv : std_logic_vector(1650 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1651_t(x : std_logic_vector) return int1651_t is
  variable rv : int1651_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1652_t_to_slv(x : uint1652_t) return std_logic_vector is
  variable rv : std_logic_vector(1651 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1652_t(x : std_logic_vector) return uint1652_t is
  variable rv : uint1652_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1652_t_to_slv(x : int1652_t) return std_logic_vector is
  variable rv : std_logic_vector(1651 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1652_t(x : std_logic_vector) return int1652_t is
  variable rv : int1652_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1653_t_to_slv(x : uint1653_t) return std_logic_vector is
  variable rv : std_logic_vector(1652 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1653_t(x : std_logic_vector) return uint1653_t is
  variable rv : uint1653_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1653_t_to_slv(x : int1653_t) return std_logic_vector is
  variable rv : std_logic_vector(1652 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1653_t(x : std_logic_vector) return int1653_t is
  variable rv : int1653_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1654_t_to_slv(x : uint1654_t) return std_logic_vector is
  variable rv : std_logic_vector(1653 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1654_t(x : std_logic_vector) return uint1654_t is
  variable rv : uint1654_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1654_t_to_slv(x : int1654_t) return std_logic_vector is
  variable rv : std_logic_vector(1653 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1654_t(x : std_logic_vector) return int1654_t is
  variable rv : int1654_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1655_t_to_slv(x : uint1655_t) return std_logic_vector is
  variable rv : std_logic_vector(1654 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1655_t(x : std_logic_vector) return uint1655_t is
  variable rv : uint1655_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1655_t_to_slv(x : int1655_t) return std_logic_vector is
  variable rv : std_logic_vector(1654 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1655_t(x : std_logic_vector) return int1655_t is
  variable rv : int1655_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1656_t_to_slv(x : uint1656_t) return std_logic_vector is
  variable rv : std_logic_vector(1655 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1656_t(x : std_logic_vector) return uint1656_t is
  variable rv : uint1656_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1656_t_to_slv(x : int1656_t) return std_logic_vector is
  variable rv : std_logic_vector(1655 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1656_t(x : std_logic_vector) return int1656_t is
  variable rv : int1656_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1657_t_to_slv(x : uint1657_t) return std_logic_vector is
  variable rv : std_logic_vector(1656 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1657_t(x : std_logic_vector) return uint1657_t is
  variable rv : uint1657_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1657_t_to_slv(x : int1657_t) return std_logic_vector is
  variable rv : std_logic_vector(1656 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1657_t(x : std_logic_vector) return int1657_t is
  variable rv : int1657_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1658_t_to_slv(x : uint1658_t) return std_logic_vector is
  variable rv : std_logic_vector(1657 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1658_t(x : std_logic_vector) return uint1658_t is
  variable rv : uint1658_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1658_t_to_slv(x : int1658_t) return std_logic_vector is
  variable rv : std_logic_vector(1657 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1658_t(x : std_logic_vector) return int1658_t is
  variable rv : int1658_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1659_t_to_slv(x : uint1659_t) return std_logic_vector is
  variable rv : std_logic_vector(1658 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1659_t(x : std_logic_vector) return uint1659_t is
  variable rv : uint1659_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1659_t_to_slv(x : int1659_t) return std_logic_vector is
  variable rv : std_logic_vector(1658 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1659_t(x : std_logic_vector) return int1659_t is
  variable rv : int1659_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1660_t_to_slv(x : uint1660_t) return std_logic_vector is
  variable rv : std_logic_vector(1659 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1660_t(x : std_logic_vector) return uint1660_t is
  variable rv : uint1660_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1660_t_to_slv(x : int1660_t) return std_logic_vector is
  variable rv : std_logic_vector(1659 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1660_t(x : std_logic_vector) return int1660_t is
  variable rv : int1660_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1661_t_to_slv(x : uint1661_t) return std_logic_vector is
  variable rv : std_logic_vector(1660 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1661_t(x : std_logic_vector) return uint1661_t is
  variable rv : uint1661_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1661_t_to_slv(x : int1661_t) return std_logic_vector is
  variable rv : std_logic_vector(1660 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1661_t(x : std_logic_vector) return int1661_t is
  variable rv : int1661_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1662_t_to_slv(x : uint1662_t) return std_logic_vector is
  variable rv : std_logic_vector(1661 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1662_t(x : std_logic_vector) return uint1662_t is
  variable rv : uint1662_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1662_t_to_slv(x : int1662_t) return std_logic_vector is
  variable rv : std_logic_vector(1661 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1662_t(x : std_logic_vector) return int1662_t is
  variable rv : int1662_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1663_t_to_slv(x : uint1663_t) return std_logic_vector is
  variable rv : std_logic_vector(1662 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1663_t(x : std_logic_vector) return uint1663_t is
  variable rv : uint1663_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1663_t_to_slv(x : int1663_t) return std_logic_vector is
  variable rv : std_logic_vector(1662 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1663_t(x : std_logic_vector) return int1663_t is
  variable rv : int1663_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1664_t_to_slv(x : uint1664_t) return std_logic_vector is
  variable rv : std_logic_vector(1663 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1664_t(x : std_logic_vector) return uint1664_t is
  variable rv : uint1664_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1664_t_to_slv(x : int1664_t) return std_logic_vector is
  variable rv : std_logic_vector(1663 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1664_t(x : std_logic_vector) return int1664_t is
  variable rv : int1664_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1665_t_to_slv(x : uint1665_t) return std_logic_vector is
  variable rv : std_logic_vector(1664 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1665_t(x : std_logic_vector) return uint1665_t is
  variable rv : uint1665_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1665_t_to_slv(x : int1665_t) return std_logic_vector is
  variable rv : std_logic_vector(1664 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1665_t(x : std_logic_vector) return int1665_t is
  variable rv : int1665_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1666_t_to_slv(x : uint1666_t) return std_logic_vector is
  variable rv : std_logic_vector(1665 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1666_t(x : std_logic_vector) return uint1666_t is
  variable rv : uint1666_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1666_t_to_slv(x : int1666_t) return std_logic_vector is
  variable rv : std_logic_vector(1665 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1666_t(x : std_logic_vector) return int1666_t is
  variable rv : int1666_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1667_t_to_slv(x : uint1667_t) return std_logic_vector is
  variable rv : std_logic_vector(1666 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1667_t(x : std_logic_vector) return uint1667_t is
  variable rv : uint1667_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1667_t_to_slv(x : int1667_t) return std_logic_vector is
  variable rv : std_logic_vector(1666 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1667_t(x : std_logic_vector) return int1667_t is
  variable rv : int1667_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1668_t_to_slv(x : uint1668_t) return std_logic_vector is
  variable rv : std_logic_vector(1667 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1668_t(x : std_logic_vector) return uint1668_t is
  variable rv : uint1668_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1668_t_to_slv(x : int1668_t) return std_logic_vector is
  variable rv : std_logic_vector(1667 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1668_t(x : std_logic_vector) return int1668_t is
  variable rv : int1668_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1669_t_to_slv(x : uint1669_t) return std_logic_vector is
  variable rv : std_logic_vector(1668 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1669_t(x : std_logic_vector) return uint1669_t is
  variable rv : uint1669_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1669_t_to_slv(x : int1669_t) return std_logic_vector is
  variable rv : std_logic_vector(1668 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1669_t(x : std_logic_vector) return int1669_t is
  variable rv : int1669_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1670_t_to_slv(x : uint1670_t) return std_logic_vector is
  variable rv : std_logic_vector(1669 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1670_t(x : std_logic_vector) return uint1670_t is
  variable rv : uint1670_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1670_t_to_slv(x : int1670_t) return std_logic_vector is
  variable rv : std_logic_vector(1669 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1670_t(x : std_logic_vector) return int1670_t is
  variable rv : int1670_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1671_t_to_slv(x : uint1671_t) return std_logic_vector is
  variable rv : std_logic_vector(1670 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1671_t(x : std_logic_vector) return uint1671_t is
  variable rv : uint1671_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1671_t_to_slv(x : int1671_t) return std_logic_vector is
  variable rv : std_logic_vector(1670 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1671_t(x : std_logic_vector) return int1671_t is
  variable rv : int1671_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1672_t_to_slv(x : uint1672_t) return std_logic_vector is
  variable rv : std_logic_vector(1671 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1672_t(x : std_logic_vector) return uint1672_t is
  variable rv : uint1672_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1672_t_to_slv(x : int1672_t) return std_logic_vector is
  variable rv : std_logic_vector(1671 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1672_t(x : std_logic_vector) return int1672_t is
  variable rv : int1672_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1673_t_to_slv(x : uint1673_t) return std_logic_vector is
  variable rv : std_logic_vector(1672 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1673_t(x : std_logic_vector) return uint1673_t is
  variable rv : uint1673_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1673_t_to_slv(x : int1673_t) return std_logic_vector is
  variable rv : std_logic_vector(1672 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1673_t(x : std_logic_vector) return int1673_t is
  variable rv : int1673_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1674_t_to_slv(x : uint1674_t) return std_logic_vector is
  variable rv : std_logic_vector(1673 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1674_t(x : std_logic_vector) return uint1674_t is
  variable rv : uint1674_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1674_t_to_slv(x : int1674_t) return std_logic_vector is
  variable rv : std_logic_vector(1673 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1674_t(x : std_logic_vector) return int1674_t is
  variable rv : int1674_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1675_t_to_slv(x : uint1675_t) return std_logic_vector is
  variable rv : std_logic_vector(1674 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1675_t(x : std_logic_vector) return uint1675_t is
  variable rv : uint1675_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1675_t_to_slv(x : int1675_t) return std_logic_vector is
  variable rv : std_logic_vector(1674 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1675_t(x : std_logic_vector) return int1675_t is
  variable rv : int1675_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1676_t_to_slv(x : uint1676_t) return std_logic_vector is
  variable rv : std_logic_vector(1675 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1676_t(x : std_logic_vector) return uint1676_t is
  variable rv : uint1676_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1676_t_to_slv(x : int1676_t) return std_logic_vector is
  variable rv : std_logic_vector(1675 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1676_t(x : std_logic_vector) return int1676_t is
  variable rv : int1676_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1677_t_to_slv(x : uint1677_t) return std_logic_vector is
  variable rv : std_logic_vector(1676 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1677_t(x : std_logic_vector) return uint1677_t is
  variable rv : uint1677_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1677_t_to_slv(x : int1677_t) return std_logic_vector is
  variable rv : std_logic_vector(1676 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1677_t(x : std_logic_vector) return int1677_t is
  variable rv : int1677_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1678_t_to_slv(x : uint1678_t) return std_logic_vector is
  variable rv : std_logic_vector(1677 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1678_t(x : std_logic_vector) return uint1678_t is
  variable rv : uint1678_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1678_t_to_slv(x : int1678_t) return std_logic_vector is
  variable rv : std_logic_vector(1677 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1678_t(x : std_logic_vector) return int1678_t is
  variable rv : int1678_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1679_t_to_slv(x : uint1679_t) return std_logic_vector is
  variable rv : std_logic_vector(1678 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1679_t(x : std_logic_vector) return uint1679_t is
  variable rv : uint1679_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1679_t_to_slv(x : int1679_t) return std_logic_vector is
  variable rv : std_logic_vector(1678 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1679_t(x : std_logic_vector) return int1679_t is
  variable rv : int1679_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1680_t_to_slv(x : uint1680_t) return std_logic_vector is
  variable rv : std_logic_vector(1679 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1680_t(x : std_logic_vector) return uint1680_t is
  variable rv : uint1680_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1680_t_to_slv(x : int1680_t) return std_logic_vector is
  variable rv : std_logic_vector(1679 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1680_t(x : std_logic_vector) return int1680_t is
  variable rv : int1680_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1681_t_to_slv(x : uint1681_t) return std_logic_vector is
  variable rv : std_logic_vector(1680 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1681_t(x : std_logic_vector) return uint1681_t is
  variable rv : uint1681_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1681_t_to_slv(x : int1681_t) return std_logic_vector is
  variable rv : std_logic_vector(1680 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1681_t(x : std_logic_vector) return int1681_t is
  variable rv : int1681_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1682_t_to_slv(x : uint1682_t) return std_logic_vector is
  variable rv : std_logic_vector(1681 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1682_t(x : std_logic_vector) return uint1682_t is
  variable rv : uint1682_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1682_t_to_slv(x : int1682_t) return std_logic_vector is
  variable rv : std_logic_vector(1681 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1682_t(x : std_logic_vector) return int1682_t is
  variable rv : int1682_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1683_t_to_slv(x : uint1683_t) return std_logic_vector is
  variable rv : std_logic_vector(1682 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1683_t(x : std_logic_vector) return uint1683_t is
  variable rv : uint1683_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1683_t_to_slv(x : int1683_t) return std_logic_vector is
  variable rv : std_logic_vector(1682 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1683_t(x : std_logic_vector) return int1683_t is
  variable rv : int1683_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1684_t_to_slv(x : uint1684_t) return std_logic_vector is
  variable rv : std_logic_vector(1683 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1684_t(x : std_logic_vector) return uint1684_t is
  variable rv : uint1684_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1684_t_to_slv(x : int1684_t) return std_logic_vector is
  variable rv : std_logic_vector(1683 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1684_t(x : std_logic_vector) return int1684_t is
  variable rv : int1684_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1685_t_to_slv(x : uint1685_t) return std_logic_vector is
  variable rv : std_logic_vector(1684 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1685_t(x : std_logic_vector) return uint1685_t is
  variable rv : uint1685_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1685_t_to_slv(x : int1685_t) return std_logic_vector is
  variable rv : std_logic_vector(1684 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1685_t(x : std_logic_vector) return int1685_t is
  variable rv : int1685_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1686_t_to_slv(x : uint1686_t) return std_logic_vector is
  variable rv : std_logic_vector(1685 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1686_t(x : std_logic_vector) return uint1686_t is
  variable rv : uint1686_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1686_t_to_slv(x : int1686_t) return std_logic_vector is
  variable rv : std_logic_vector(1685 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1686_t(x : std_logic_vector) return int1686_t is
  variable rv : int1686_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1687_t_to_slv(x : uint1687_t) return std_logic_vector is
  variable rv : std_logic_vector(1686 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1687_t(x : std_logic_vector) return uint1687_t is
  variable rv : uint1687_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1687_t_to_slv(x : int1687_t) return std_logic_vector is
  variable rv : std_logic_vector(1686 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1687_t(x : std_logic_vector) return int1687_t is
  variable rv : int1687_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1688_t_to_slv(x : uint1688_t) return std_logic_vector is
  variable rv : std_logic_vector(1687 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1688_t(x : std_logic_vector) return uint1688_t is
  variable rv : uint1688_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1688_t_to_slv(x : int1688_t) return std_logic_vector is
  variable rv : std_logic_vector(1687 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1688_t(x : std_logic_vector) return int1688_t is
  variable rv : int1688_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1689_t_to_slv(x : uint1689_t) return std_logic_vector is
  variable rv : std_logic_vector(1688 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1689_t(x : std_logic_vector) return uint1689_t is
  variable rv : uint1689_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1689_t_to_slv(x : int1689_t) return std_logic_vector is
  variable rv : std_logic_vector(1688 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1689_t(x : std_logic_vector) return int1689_t is
  variable rv : int1689_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1690_t_to_slv(x : uint1690_t) return std_logic_vector is
  variable rv : std_logic_vector(1689 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1690_t(x : std_logic_vector) return uint1690_t is
  variable rv : uint1690_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1690_t_to_slv(x : int1690_t) return std_logic_vector is
  variable rv : std_logic_vector(1689 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1690_t(x : std_logic_vector) return int1690_t is
  variable rv : int1690_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1691_t_to_slv(x : uint1691_t) return std_logic_vector is
  variable rv : std_logic_vector(1690 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1691_t(x : std_logic_vector) return uint1691_t is
  variable rv : uint1691_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1691_t_to_slv(x : int1691_t) return std_logic_vector is
  variable rv : std_logic_vector(1690 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1691_t(x : std_logic_vector) return int1691_t is
  variable rv : int1691_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1692_t_to_slv(x : uint1692_t) return std_logic_vector is
  variable rv : std_logic_vector(1691 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1692_t(x : std_logic_vector) return uint1692_t is
  variable rv : uint1692_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1692_t_to_slv(x : int1692_t) return std_logic_vector is
  variable rv : std_logic_vector(1691 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1692_t(x : std_logic_vector) return int1692_t is
  variable rv : int1692_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1693_t_to_slv(x : uint1693_t) return std_logic_vector is
  variable rv : std_logic_vector(1692 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1693_t(x : std_logic_vector) return uint1693_t is
  variable rv : uint1693_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1693_t_to_slv(x : int1693_t) return std_logic_vector is
  variable rv : std_logic_vector(1692 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1693_t(x : std_logic_vector) return int1693_t is
  variable rv : int1693_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1694_t_to_slv(x : uint1694_t) return std_logic_vector is
  variable rv : std_logic_vector(1693 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1694_t(x : std_logic_vector) return uint1694_t is
  variable rv : uint1694_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1694_t_to_slv(x : int1694_t) return std_logic_vector is
  variable rv : std_logic_vector(1693 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1694_t(x : std_logic_vector) return int1694_t is
  variable rv : int1694_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1695_t_to_slv(x : uint1695_t) return std_logic_vector is
  variable rv : std_logic_vector(1694 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1695_t(x : std_logic_vector) return uint1695_t is
  variable rv : uint1695_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1695_t_to_slv(x : int1695_t) return std_logic_vector is
  variable rv : std_logic_vector(1694 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1695_t(x : std_logic_vector) return int1695_t is
  variable rv : int1695_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1696_t_to_slv(x : uint1696_t) return std_logic_vector is
  variable rv : std_logic_vector(1695 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1696_t(x : std_logic_vector) return uint1696_t is
  variable rv : uint1696_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1696_t_to_slv(x : int1696_t) return std_logic_vector is
  variable rv : std_logic_vector(1695 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1696_t(x : std_logic_vector) return int1696_t is
  variable rv : int1696_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1697_t_to_slv(x : uint1697_t) return std_logic_vector is
  variable rv : std_logic_vector(1696 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1697_t(x : std_logic_vector) return uint1697_t is
  variable rv : uint1697_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1697_t_to_slv(x : int1697_t) return std_logic_vector is
  variable rv : std_logic_vector(1696 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1697_t(x : std_logic_vector) return int1697_t is
  variable rv : int1697_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1698_t_to_slv(x : uint1698_t) return std_logic_vector is
  variable rv : std_logic_vector(1697 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1698_t(x : std_logic_vector) return uint1698_t is
  variable rv : uint1698_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1698_t_to_slv(x : int1698_t) return std_logic_vector is
  variable rv : std_logic_vector(1697 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1698_t(x : std_logic_vector) return int1698_t is
  variable rv : int1698_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1699_t_to_slv(x : uint1699_t) return std_logic_vector is
  variable rv : std_logic_vector(1698 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1699_t(x : std_logic_vector) return uint1699_t is
  variable rv : uint1699_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1699_t_to_slv(x : int1699_t) return std_logic_vector is
  variable rv : std_logic_vector(1698 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1699_t(x : std_logic_vector) return int1699_t is
  variable rv : int1699_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1700_t_to_slv(x : uint1700_t) return std_logic_vector is
  variable rv : std_logic_vector(1699 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1700_t(x : std_logic_vector) return uint1700_t is
  variable rv : uint1700_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1700_t_to_slv(x : int1700_t) return std_logic_vector is
  variable rv : std_logic_vector(1699 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1700_t(x : std_logic_vector) return int1700_t is
  variable rv : int1700_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1701_t_to_slv(x : uint1701_t) return std_logic_vector is
  variable rv : std_logic_vector(1700 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1701_t(x : std_logic_vector) return uint1701_t is
  variable rv : uint1701_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1701_t_to_slv(x : int1701_t) return std_logic_vector is
  variable rv : std_logic_vector(1700 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1701_t(x : std_logic_vector) return int1701_t is
  variable rv : int1701_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1702_t_to_slv(x : uint1702_t) return std_logic_vector is
  variable rv : std_logic_vector(1701 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1702_t(x : std_logic_vector) return uint1702_t is
  variable rv : uint1702_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1702_t_to_slv(x : int1702_t) return std_logic_vector is
  variable rv : std_logic_vector(1701 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1702_t(x : std_logic_vector) return int1702_t is
  variable rv : int1702_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1703_t_to_slv(x : uint1703_t) return std_logic_vector is
  variable rv : std_logic_vector(1702 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1703_t(x : std_logic_vector) return uint1703_t is
  variable rv : uint1703_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1703_t_to_slv(x : int1703_t) return std_logic_vector is
  variable rv : std_logic_vector(1702 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1703_t(x : std_logic_vector) return int1703_t is
  variable rv : int1703_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1704_t_to_slv(x : uint1704_t) return std_logic_vector is
  variable rv : std_logic_vector(1703 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1704_t(x : std_logic_vector) return uint1704_t is
  variable rv : uint1704_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1704_t_to_slv(x : int1704_t) return std_logic_vector is
  variable rv : std_logic_vector(1703 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1704_t(x : std_logic_vector) return int1704_t is
  variable rv : int1704_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1705_t_to_slv(x : uint1705_t) return std_logic_vector is
  variable rv : std_logic_vector(1704 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1705_t(x : std_logic_vector) return uint1705_t is
  variable rv : uint1705_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1705_t_to_slv(x : int1705_t) return std_logic_vector is
  variable rv : std_logic_vector(1704 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1705_t(x : std_logic_vector) return int1705_t is
  variable rv : int1705_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1706_t_to_slv(x : uint1706_t) return std_logic_vector is
  variable rv : std_logic_vector(1705 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1706_t(x : std_logic_vector) return uint1706_t is
  variable rv : uint1706_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1706_t_to_slv(x : int1706_t) return std_logic_vector is
  variable rv : std_logic_vector(1705 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1706_t(x : std_logic_vector) return int1706_t is
  variable rv : int1706_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1707_t_to_slv(x : uint1707_t) return std_logic_vector is
  variable rv : std_logic_vector(1706 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1707_t(x : std_logic_vector) return uint1707_t is
  variable rv : uint1707_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1707_t_to_slv(x : int1707_t) return std_logic_vector is
  variable rv : std_logic_vector(1706 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1707_t(x : std_logic_vector) return int1707_t is
  variable rv : int1707_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1708_t_to_slv(x : uint1708_t) return std_logic_vector is
  variable rv : std_logic_vector(1707 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1708_t(x : std_logic_vector) return uint1708_t is
  variable rv : uint1708_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1708_t_to_slv(x : int1708_t) return std_logic_vector is
  variable rv : std_logic_vector(1707 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1708_t(x : std_logic_vector) return int1708_t is
  variable rv : int1708_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1709_t_to_slv(x : uint1709_t) return std_logic_vector is
  variable rv : std_logic_vector(1708 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1709_t(x : std_logic_vector) return uint1709_t is
  variable rv : uint1709_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1709_t_to_slv(x : int1709_t) return std_logic_vector is
  variable rv : std_logic_vector(1708 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1709_t(x : std_logic_vector) return int1709_t is
  variable rv : int1709_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1710_t_to_slv(x : uint1710_t) return std_logic_vector is
  variable rv : std_logic_vector(1709 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1710_t(x : std_logic_vector) return uint1710_t is
  variable rv : uint1710_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1710_t_to_slv(x : int1710_t) return std_logic_vector is
  variable rv : std_logic_vector(1709 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1710_t(x : std_logic_vector) return int1710_t is
  variable rv : int1710_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1711_t_to_slv(x : uint1711_t) return std_logic_vector is
  variable rv : std_logic_vector(1710 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1711_t(x : std_logic_vector) return uint1711_t is
  variable rv : uint1711_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1711_t_to_slv(x : int1711_t) return std_logic_vector is
  variable rv : std_logic_vector(1710 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1711_t(x : std_logic_vector) return int1711_t is
  variable rv : int1711_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1712_t_to_slv(x : uint1712_t) return std_logic_vector is
  variable rv : std_logic_vector(1711 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1712_t(x : std_logic_vector) return uint1712_t is
  variable rv : uint1712_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1712_t_to_slv(x : int1712_t) return std_logic_vector is
  variable rv : std_logic_vector(1711 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1712_t(x : std_logic_vector) return int1712_t is
  variable rv : int1712_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1713_t_to_slv(x : uint1713_t) return std_logic_vector is
  variable rv : std_logic_vector(1712 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1713_t(x : std_logic_vector) return uint1713_t is
  variable rv : uint1713_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1713_t_to_slv(x : int1713_t) return std_logic_vector is
  variable rv : std_logic_vector(1712 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1713_t(x : std_logic_vector) return int1713_t is
  variable rv : int1713_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1714_t_to_slv(x : uint1714_t) return std_logic_vector is
  variable rv : std_logic_vector(1713 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1714_t(x : std_logic_vector) return uint1714_t is
  variable rv : uint1714_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1714_t_to_slv(x : int1714_t) return std_logic_vector is
  variable rv : std_logic_vector(1713 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1714_t(x : std_logic_vector) return int1714_t is
  variable rv : int1714_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1715_t_to_slv(x : uint1715_t) return std_logic_vector is
  variable rv : std_logic_vector(1714 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1715_t(x : std_logic_vector) return uint1715_t is
  variable rv : uint1715_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1715_t_to_slv(x : int1715_t) return std_logic_vector is
  variable rv : std_logic_vector(1714 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1715_t(x : std_logic_vector) return int1715_t is
  variable rv : int1715_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1716_t_to_slv(x : uint1716_t) return std_logic_vector is
  variable rv : std_logic_vector(1715 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1716_t(x : std_logic_vector) return uint1716_t is
  variable rv : uint1716_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1716_t_to_slv(x : int1716_t) return std_logic_vector is
  variable rv : std_logic_vector(1715 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1716_t(x : std_logic_vector) return int1716_t is
  variable rv : int1716_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1717_t_to_slv(x : uint1717_t) return std_logic_vector is
  variable rv : std_logic_vector(1716 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1717_t(x : std_logic_vector) return uint1717_t is
  variable rv : uint1717_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1717_t_to_slv(x : int1717_t) return std_logic_vector is
  variable rv : std_logic_vector(1716 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1717_t(x : std_logic_vector) return int1717_t is
  variable rv : int1717_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1718_t_to_slv(x : uint1718_t) return std_logic_vector is
  variable rv : std_logic_vector(1717 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1718_t(x : std_logic_vector) return uint1718_t is
  variable rv : uint1718_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1718_t_to_slv(x : int1718_t) return std_logic_vector is
  variable rv : std_logic_vector(1717 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1718_t(x : std_logic_vector) return int1718_t is
  variable rv : int1718_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1719_t_to_slv(x : uint1719_t) return std_logic_vector is
  variable rv : std_logic_vector(1718 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1719_t(x : std_logic_vector) return uint1719_t is
  variable rv : uint1719_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1719_t_to_slv(x : int1719_t) return std_logic_vector is
  variable rv : std_logic_vector(1718 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1719_t(x : std_logic_vector) return int1719_t is
  variable rv : int1719_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1720_t_to_slv(x : uint1720_t) return std_logic_vector is
  variable rv : std_logic_vector(1719 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1720_t(x : std_logic_vector) return uint1720_t is
  variable rv : uint1720_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1720_t_to_slv(x : int1720_t) return std_logic_vector is
  variable rv : std_logic_vector(1719 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1720_t(x : std_logic_vector) return int1720_t is
  variable rv : int1720_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1721_t_to_slv(x : uint1721_t) return std_logic_vector is
  variable rv : std_logic_vector(1720 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1721_t(x : std_logic_vector) return uint1721_t is
  variable rv : uint1721_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1721_t_to_slv(x : int1721_t) return std_logic_vector is
  variable rv : std_logic_vector(1720 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1721_t(x : std_logic_vector) return int1721_t is
  variable rv : int1721_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1722_t_to_slv(x : uint1722_t) return std_logic_vector is
  variable rv : std_logic_vector(1721 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1722_t(x : std_logic_vector) return uint1722_t is
  variable rv : uint1722_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1722_t_to_slv(x : int1722_t) return std_logic_vector is
  variable rv : std_logic_vector(1721 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1722_t(x : std_logic_vector) return int1722_t is
  variable rv : int1722_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1723_t_to_slv(x : uint1723_t) return std_logic_vector is
  variable rv : std_logic_vector(1722 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1723_t(x : std_logic_vector) return uint1723_t is
  variable rv : uint1723_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1723_t_to_slv(x : int1723_t) return std_logic_vector is
  variable rv : std_logic_vector(1722 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1723_t(x : std_logic_vector) return int1723_t is
  variable rv : int1723_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1724_t_to_slv(x : uint1724_t) return std_logic_vector is
  variable rv : std_logic_vector(1723 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1724_t(x : std_logic_vector) return uint1724_t is
  variable rv : uint1724_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1724_t_to_slv(x : int1724_t) return std_logic_vector is
  variable rv : std_logic_vector(1723 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1724_t(x : std_logic_vector) return int1724_t is
  variable rv : int1724_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1725_t_to_slv(x : uint1725_t) return std_logic_vector is
  variable rv : std_logic_vector(1724 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1725_t(x : std_logic_vector) return uint1725_t is
  variable rv : uint1725_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1725_t_to_slv(x : int1725_t) return std_logic_vector is
  variable rv : std_logic_vector(1724 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1725_t(x : std_logic_vector) return int1725_t is
  variable rv : int1725_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1726_t_to_slv(x : uint1726_t) return std_logic_vector is
  variable rv : std_logic_vector(1725 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1726_t(x : std_logic_vector) return uint1726_t is
  variable rv : uint1726_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1726_t_to_slv(x : int1726_t) return std_logic_vector is
  variable rv : std_logic_vector(1725 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1726_t(x : std_logic_vector) return int1726_t is
  variable rv : int1726_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1727_t_to_slv(x : uint1727_t) return std_logic_vector is
  variable rv : std_logic_vector(1726 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1727_t(x : std_logic_vector) return uint1727_t is
  variable rv : uint1727_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1727_t_to_slv(x : int1727_t) return std_logic_vector is
  variable rv : std_logic_vector(1726 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1727_t(x : std_logic_vector) return int1727_t is
  variable rv : int1727_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1728_t_to_slv(x : uint1728_t) return std_logic_vector is
  variable rv : std_logic_vector(1727 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1728_t(x : std_logic_vector) return uint1728_t is
  variable rv : uint1728_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1728_t_to_slv(x : int1728_t) return std_logic_vector is
  variable rv : std_logic_vector(1727 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1728_t(x : std_logic_vector) return int1728_t is
  variable rv : int1728_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1729_t_to_slv(x : uint1729_t) return std_logic_vector is
  variable rv : std_logic_vector(1728 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1729_t(x : std_logic_vector) return uint1729_t is
  variable rv : uint1729_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1729_t_to_slv(x : int1729_t) return std_logic_vector is
  variable rv : std_logic_vector(1728 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1729_t(x : std_logic_vector) return int1729_t is
  variable rv : int1729_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1730_t_to_slv(x : uint1730_t) return std_logic_vector is
  variable rv : std_logic_vector(1729 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1730_t(x : std_logic_vector) return uint1730_t is
  variable rv : uint1730_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1730_t_to_slv(x : int1730_t) return std_logic_vector is
  variable rv : std_logic_vector(1729 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1730_t(x : std_logic_vector) return int1730_t is
  variable rv : int1730_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1731_t_to_slv(x : uint1731_t) return std_logic_vector is
  variable rv : std_logic_vector(1730 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1731_t(x : std_logic_vector) return uint1731_t is
  variable rv : uint1731_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1731_t_to_slv(x : int1731_t) return std_logic_vector is
  variable rv : std_logic_vector(1730 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1731_t(x : std_logic_vector) return int1731_t is
  variable rv : int1731_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1732_t_to_slv(x : uint1732_t) return std_logic_vector is
  variable rv : std_logic_vector(1731 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1732_t(x : std_logic_vector) return uint1732_t is
  variable rv : uint1732_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1732_t_to_slv(x : int1732_t) return std_logic_vector is
  variable rv : std_logic_vector(1731 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1732_t(x : std_logic_vector) return int1732_t is
  variable rv : int1732_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1733_t_to_slv(x : uint1733_t) return std_logic_vector is
  variable rv : std_logic_vector(1732 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1733_t(x : std_logic_vector) return uint1733_t is
  variable rv : uint1733_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1733_t_to_slv(x : int1733_t) return std_logic_vector is
  variable rv : std_logic_vector(1732 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1733_t(x : std_logic_vector) return int1733_t is
  variable rv : int1733_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1734_t_to_slv(x : uint1734_t) return std_logic_vector is
  variable rv : std_logic_vector(1733 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1734_t(x : std_logic_vector) return uint1734_t is
  variable rv : uint1734_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1734_t_to_slv(x : int1734_t) return std_logic_vector is
  variable rv : std_logic_vector(1733 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1734_t(x : std_logic_vector) return int1734_t is
  variable rv : int1734_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1735_t_to_slv(x : uint1735_t) return std_logic_vector is
  variable rv : std_logic_vector(1734 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1735_t(x : std_logic_vector) return uint1735_t is
  variable rv : uint1735_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1735_t_to_slv(x : int1735_t) return std_logic_vector is
  variable rv : std_logic_vector(1734 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1735_t(x : std_logic_vector) return int1735_t is
  variable rv : int1735_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1736_t_to_slv(x : uint1736_t) return std_logic_vector is
  variable rv : std_logic_vector(1735 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1736_t(x : std_logic_vector) return uint1736_t is
  variable rv : uint1736_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1736_t_to_slv(x : int1736_t) return std_logic_vector is
  variable rv : std_logic_vector(1735 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1736_t(x : std_logic_vector) return int1736_t is
  variable rv : int1736_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1737_t_to_slv(x : uint1737_t) return std_logic_vector is
  variable rv : std_logic_vector(1736 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1737_t(x : std_logic_vector) return uint1737_t is
  variable rv : uint1737_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1737_t_to_slv(x : int1737_t) return std_logic_vector is
  variable rv : std_logic_vector(1736 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1737_t(x : std_logic_vector) return int1737_t is
  variable rv : int1737_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1738_t_to_slv(x : uint1738_t) return std_logic_vector is
  variable rv : std_logic_vector(1737 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1738_t(x : std_logic_vector) return uint1738_t is
  variable rv : uint1738_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1738_t_to_slv(x : int1738_t) return std_logic_vector is
  variable rv : std_logic_vector(1737 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1738_t(x : std_logic_vector) return int1738_t is
  variable rv : int1738_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1739_t_to_slv(x : uint1739_t) return std_logic_vector is
  variable rv : std_logic_vector(1738 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1739_t(x : std_logic_vector) return uint1739_t is
  variable rv : uint1739_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1739_t_to_slv(x : int1739_t) return std_logic_vector is
  variable rv : std_logic_vector(1738 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1739_t(x : std_logic_vector) return int1739_t is
  variable rv : int1739_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1740_t_to_slv(x : uint1740_t) return std_logic_vector is
  variable rv : std_logic_vector(1739 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1740_t(x : std_logic_vector) return uint1740_t is
  variable rv : uint1740_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1740_t_to_slv(x : int1740_t) return std_logic_vector is
  variable rv : std_logic_vector(1739 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1740_t(x : std_logic_vector) return int1740_t is
  variable rv : int1740_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1741_t_to_slv(x : uint1741_t) return std_logic_vector is
  variable rv : std_logic_vector(1740 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1741_t(x : std_logic_vector) return uint1741_t is
  variable rv : uint1741_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1741_t_to_slv(x : int1741_t) return std_logic_vector is
  variable rv : std_logic_vector(1740 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1741_t(x : std_logic_vector) return int1741_t is
  variable rv : int1741_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1742_t_to_slv(x : uint1742_t) return std_logic_vector is
  variable rv : std_logic_vector(1741 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1742_t(x : std_logic_vector) return uint1742_t is
  variable rv : uint1742_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1742_t_to_slv(x : int1742_t) return std_logic_vector is
  variable rv : std_logic_vector(1741 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1742_t(x : std_logic_vector) return int1742_t is
  variable rv : int1742_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1743_t_to_slv(x : uint1743_t) return std_logic_vector is
  variable rv : std_logic_vector(1742 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1743_t(x : std_logic_vector) return uint1743_t is
  variable rv : uint1743_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1743_t_to_slv(x : int1743_t) return std_logic_vector is
  variable rv : std_logic_vector(1742 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1743_t(x : std_logic_vector) return int1743_t is
  variable rv : int1743_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1744_t_to_slv(x : uint1744_t) return std_logic_vector is
  variable rv : std_logic_vector(1743 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1744_t(x : std_logic_vector) return uint1744_t is
  variable rv : uint1744_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1744_t_to_slv(x : int1744_t) return std_logic_vector is
  variable rv : std_logic_vector(1743 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1744_t(x : std_logic_vector) return int1744_t is
  variable rv : int1744_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1745_t_to_slv(x : uint1745_t) return std_logic_vector is
  variable rv : std_logic_vector(1744 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1745_t(x : std_logic_vector) return uint1745_t is
  variable rv : uint1745_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1745_t_to_slv(x : int1745_t) return std_logic_vector is
  variable rv : std_logic_vector(1744 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1745_t(x : std_logic_vector) return int1745_t is
  variable rv : int1745_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1746_t_to_slv(x : uint1746_t) return std_logic_vector is
  variable rv : std_logic_vector(1745 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1746_t(x : std_logic_vector) return uint1746_t is
  variable rv : uint1746_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1746_t_to_slv(x : int1746_t) return std_logic_vector is
  variable rv : std_logic_vector(1745 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1746_t(x : std_logic_vector) return int1746_t is
  variable rv : int1746_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1747_t_to_slv(x : uint1747_t) return std_logic_vector is
  variable rv : std_logic_vector(1746 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1747_t(x : std_logic_vector) return uint1747_t is
  variable rv : uint1747_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1747_t_to_slv(x : int1747_t) return std_logic_vector is
  variable rv : std_logic_vector(1746 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1747_t(x : std_logic_vector) return int1747_t is
  variable rv : int1747_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1748_t_to_slv(x : uint1748_t) return std_logic_vector is
  variable rv : std_logic_vector(1747 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1748_t(x : std_logic_vector) return uint1748_t is
  variable rv : uint1748_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1748_t_to_slv(x : int1748_t) return std_logic_vector is
  variable rv : std_logic_vector(1747 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1748_t(x : std_logic_vector) return int1748_t is
  variable rv : int1748_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1749_t_to_slv(x : uint1749_t) return std_logic_vector is
  variable rv : std_logic_vector(1748 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1749_t(x : std_logic_vector) return uint1749_t is
  variable rv : uint1749_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1749_t_to_slv(x : int1749_t) return std_logic_vector is
  variable rv : std_logic_vector(1748 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1749_t(x : std_logic_vector) return int1749_t is
  variable rv : int1749_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1750_t_to_slv(x : uint1750_t) return std_logic_vector is
  variable rv : std_logic_vector(1749 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1750_t(x : std_logic_vector) return uint1750_t is
  variable rv : uint1750_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1750_t_to_slv(x : int1750_t) return std_logic_vector is
  variable rv : std_logic_vector(1749 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1750_t(x : std_logic_vector) return int1750_t is
  variable rv : int1750_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1751_t_to_slv(x : uint1751_t) return std_logic_vector is
  variable rv : std_logic_vector(1750 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1751_t(x : std_logic_vector) return uint1751_t is
  variable rv : uint1751_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1751_t_to_slv(x : int1751_t) return std_logic_vector is
  variable rv : std_logic_vector(1750 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1751_t(x : std_logic_vector) return int1751_t is
  variable rv : int1751_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1752_t_to_slv(x : uint1752_t) return std_logic_vector is
  variable rv : std_logic_vector(1751 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1752_t(x : std_logic_vector) return uint1752_t is
  variable rv : uint1752_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1752_t_to_slv(x : int1752_t) return std_logic_vector is
  variable rv : std_logic_vector(1751 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1752_t(x : std_logic_vector) return int1752_t is
  variable rv : int1752_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1753_t_to_slv(x : uint1753_t) return std_logic_vector is
  variable rv : std_logic_vector(1752 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1753_t(x : std_logic_vector) return uint1753_t is
  variable rv : uint1753_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1753_t_to_slv(x : int1753_t) return std_logic_vector is
  variable rv : std_logic_vector(1752 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1753_t(x : std_logic_vector) return int1753_t is
  variable rv : int1753_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1754_t_to_slv(x : uint1754_t) return std_logic_vector is
  variable rv : std_logic_vector(1753 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1754_t(x : std_logic_vector) return uint1754_t is
  variable rv : uint1754_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1754_t_to_slv(x : int1754_t) return std_logic_vector is
  variable rv : std_logic_vector(1753 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1754_t(x : std_logic_vector) return int1754_t is
  variable rv : int1754_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1755_t_to_slv(x : uint1755_t) return std_logic_vector is
  variable rv : std_logic_vector(1754 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1755_t(x : std_logic_vector) return uint1755_t is
  variable rv : uint1755_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1755_t_to_slv(x : int1755_t) return std_logic_vector is
  variable rv : std_logic_vector(1754 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1755_t(x : std_logic_vector) return int1755_t is
  variable rv : int1755_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1756_t_to_slv(x : uint1756_t) return std_logic_vector is
  variable rv : std_logic_vector(1755 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1756_t(x : std_logic_vector) return uint1756_t is
  variable rv : uint1756_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1756_t_to_slv(x : int1756_t) return std_logic_vector is
  variable rv : std_logic_vector(1755 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1756_t(x : std_logic_vector) return int1756_t is
  variable rv : int1756_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1757_t_to_slv(x : uint1757_t) return std_logic_vector is
  variable rv : std_logic_vector(1756 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1757_t(x : std_logic_vector) return uint1757_t is
  variable rv : uint1757_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1757_t_to_slv(x : int1757_t) return std_logic_vector is
  variable rv : std_logic_vector(1756 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1757_t(x : std_logic_vector) return int1757_t is
  variable rv : int1757_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1758_t_to_slv(x : uint1758_t) return std_logic_vector is
  variable rv : std_logic_vector(1757 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1758_t(x : std_logic_vector) return uint1758_t is
  variable rv : uint1758_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1758_t_to_slv(x : int1758_t) return std_logic_vector is
  variable rv : std_logic_vector(1757 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1758_t(x : std_logic_vector) return int1758_t is
  variable rv : int1758_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1759_t_to_slv(x : uint1759_t) return std_logic_vector is
  variable rv : std_logic_vector(1758 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1759_t(x : std_logic_vector) return uint1759_t is
  variable rv : uint1759_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1759_t_to_slv(x : int1759_t) return std_logic_vector is
  variable rv : std_logic_vector(1758 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1759_t(x : std_logic_vector) return int1759_t is
  variable rv : int1759_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1760_t_to_slv(x : uint1760_t) return std_logic_vector is
  variable rv : std_logic_vector(1759 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1760_t(x : std_logic_vector) return uint1760_t is
  variable rv : uint1760_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1760_t_to_slv(x : int1760_t) return std_logic_vector is
  variable rv : std_logic_vector(1759 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1760_t(x : std_logic_vector) return int1760_t is
  variable rv : int1760_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1761_t_to_slv(x : uint1761_t) return std_logic_vector is
  variable rv : std_logic_vector(1760 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1761_t(x : std_logic_vector) return uint1761_t is
  variable rv : uint1761_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1761_t_to_slv(x : int1761_t) return std_logic_vector is
  variable rv : std_logic_vector(1760 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1761_t(x : std_logic_vector) return int1761_t is
  variable rv : int1761_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1762_t_to_slv(x : uint1762_t) return std_logic_vector is
  variable rv : std_logic_vector(1761 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1762_t(x : std_logic_vector) return uint1762_t is
  variable rv : uint1762_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1762_t_to_slv(x : int1762_t) return std_logic_vector is
  variable rv : std_logic_vector(1761 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1762_t(x : std_logic_vector) return int1762_t is
  variable rv : int1762_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1763_t_to_slv(x : uint1763_t) return std_logic_vector is
  variable rv : std_logic_vector(1762 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1763_t(x : std_logic_vector) return uint1763_t is
  variable rv : uint1763_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1763_t_to_slv(x : int1763_t) return std_logic_vector is
  variable rv : std_logic_vector(1762 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1763_t(x : std_logic_vector) return int1763_t is
  variable rv : int1763_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1764_t_to_slv(x : uint1764_t) return std_logic_vector is
  variable rv : std_logic_vector(1763 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1764_t(x : std_logic_vector) return uint1764_t is
  variable rv : uint1764_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1764_t_to_slv(x : int1764_t) return std_logic_vector is
  variable rv : std_logic_vector(1763 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1764_t(x : std_logic_vector) return int1764_t is
  variable rv : int1764_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1765_t_to_slv(x : uint1765_t) return std_logic_vector is
  variable rv : std_logic_vector(1764 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1765_t(x : std_logic_vector) return uint1765_t is
  variable rv : uint1765_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1765_t_to_slv(x : int1765_t) return std_logic_vector is
  variable rv : std_logic_vector(1764 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1765_t(x : std_logic_vector) return int1765_t is
  variable rv : int1765_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1766_t_to_slv(x : uint1766_t) return std_logic_vector is
  variable rv : std_logic_vector(1765 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1766_t(x : std_logic_vector) return uint1766_t is
  variable rv : uint1766_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1766_t_to_slv(x : int1766_t) return std_logic_vector is
  variable rv : std_logic_vector(1765 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1766_t(x : std_logic_vector) return int1766_t is
  variable rv : int1766_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1767_t_to_slv(x : uint1767_t) return std_logic_vector is
  variable rv : std_logic_vector(1766 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1767_t(x : std_logic_vector) return uint1767_t is
  variable rv : uint1767_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1767_t_to_slv(x : int1767_t) return std_logic_vector is
  variable rv : std_logic_vector(1766 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1767_t(x : std_logic_vector) return int1767_t is
  variable rv : int1767_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1768_t_to_slv(x : uint1768_t) return std_logic_vector is
  variable rv : std_logic_vector(1767 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1768_t(x : std_logic_vector) return uint1768_t is
  variable rv : uint1768_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1768_t_to_slv(x : int1768_t) return std_logic_vector is
  variable rv : std_logic_vector(1767 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1768_t(x : std_logic_vector) return int1768_t is
  variable rv : int1768_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1769_t_to_slv(x : uint1769_t) return std_logic_vector is
  variable rv : std_logic_vector(1768 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1769_t(x : std_logic_vector) return uint1769_t is
  variable rv : uint1769_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1769_t_to_slv(x : int1769_t) return std_logic_vector is
  variable rv : std_logic_vector(1768 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1769_t(x : std_logic_vector) return int1769_t is
  variable rv : int1769_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1770_t_to_slv(x : uint1770_t) return std_logic_vector is
  variable rv : std_logic_vector(1769 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1770_t(x : std_logic_vector) return uint1770_t is
  variable rv : uint1770_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1770_t_to_slv(x : int1770_t) return std_logic_vector is
  variable rv : std_logic_vector(1769 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1770_t(x : std_logic_vector) return int1770_t is
  variable rv : int1770_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1771_t_to_slv(x : uint1771_t) return std_logic_vector is
  variable rv : std_logic_vector(1770 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1771_t(x : std_logic_vector) return uint1771_t is
  variable rv : uint1771_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1771_t_to_slv(x : int1771_t) return std_logic_vector is
  variable rv : std_logic_vector(1770 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1771_t(x : std_logic_vector) return int1771_t is
  variable rv : int1771_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1772_t_to_slv(x : uint1772_t) return std_logic_vector is
  variable rv : std_logic_vector(1771 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1772_t(x : std_logic_vector) return uint1772_t is
  variable rv : uint1772_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1772_t_to_slv(x : int1772_t) return std_logic_vector is
  variable rv : std_logic_vector(1771 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1772_t(x : std_logic_vector) return int1772_t is
  variable rv : int1772_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1773_t_to_slv(x : uint1773_t) return std_logic_vector is
  variable rv : std_logic_vector(1772 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1773_t(x : std_logic_vector) return uint1773_t is
  variable rv : uint1773_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1773_t_to_slv(x : int1773_t) return std_logic_vector is
  variable rv : std_logic_vector(1772 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1773_t(x : std_logic_vector) return int1773_t is
  variable rv : int1773_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1774_t_to_slv(x : uint1774_t) return std_logic_vector is
  variable rv : std_logic_vector(1773 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1774_t(x : std_logic_vector) return uint1774_t is
  variable rv : uint1774_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1774_t_to_slv(x : int1774_t) return std_logic_vector is
  variable rv : std_logic_vector(1773 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1774_t(x : std_logic_vector) return int1774_t is
  variable rv : int1774_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1775_t_to_slv(x : uint1775_t) return std_logic_vector is
  variable rv : std_logic_vector(1774 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1775_t(x : std_logic_vector) return uint1775_t is
  variable rv : uint1775_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1775_t_to_slv(x : int1775_t) return std_logic_vector is
  variable rv : std_logic_vector(1774 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1775_t(x : std_logic_vector) return int1775_t is
  variable rv : int1775_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1776_t_to_slv(x : uint1776_t) return std_logic_vector is
  variable rv : std_logic_vector(1775 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1776_t(x : std_logic_vector) return uint1776_t is
  variable rv : uint1776_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1776_t_to_slv(x : int1776_t) return std_logic_vector is
  variable rv : std_logic_vector(1775 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1776_t(x : std_logic_vector) return int1776_t is
  variable rv : int1776_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1777_t_to_slv(x : uint1777_t) return std_logic_vector is
  variable rv : std_logic_vector(1776 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1777_t(x : std_logic_vector) return uint1777_t is
  variable rv : uint1777_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1777_t_to_slv(x : int1777_t) return std_logic_vector is
  variable rv : std_logic_vector(1776 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1777_t(x : std_logic_vector) return int1777_t is
  variable rv : int1777_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1778_t_to_slv(x : uint1778_t) return std_logic_vector is
  variable rv : std_logic_vector(1777 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1778_t(x : std_logic_vector) return uint1778_t is
  variable rv : uint1778_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1778_t_to_slv(x : int1778_t) return std_logic_vector is
  variable rv : std_logic_vector(1777 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1778_t(x : std_logic_vector) return int1778_t is
  variable rv : int1778_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1779_t_to_slv(x : uint1779_t) return std_logic_vector is
  variable rv : std_logic_vector(1778 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1779_t(x : std_logic_vector) return uint1779_t is
  variable rv : uint1779_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1779_t_to_slv(x : int1779_t) return std_logic_vector is
  variable rv : std_logic_vector(1778 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1779_t(x : std_logic_vector) return int1779_t is
  variable rv : int1779_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1780_t_to_slv(x : uint1780_t) return std_logic_vector is
  variable rv : std_logic_vector(1779 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1780_t(x : std_logic_vector) return uint1780_t is
  variable rv : uint1780_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1780_t_to_slv(x : int1780_t) return std_logic_vector is
  variable rv : std_logic_vector(1779 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1780_t(x : std_logic_vector) return int1780_t is
  variable rv : int1780_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1781_t_to_slv(x : uint1781_t) return std_logic_vector is
  variable rv : std_logic_vector(1780 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1781_t(x : std_logic_vector) return uint1781_t is
  variable rv : uint1781_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1781_t_to_slv(x : int1781_t) return std_logic_vector is
  variable rv : std_logic_vector(1780 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1781_t(x : std_logic_vector) return int1781_t is
  variable rv : int1781_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1782_t_to_slv(x : uint1782_t) return std_logic_vector is
  variable rv : std_logic_vector(1781 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1782_t(x : std_logic_vector) return uint1782_t is
  variable rv : uint1782_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1782_t_to_slv(x : int1782_t) return std_logic_vector is
  variable rv : std_logic_vector(1781 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1782_t(x : std_logic_vector) return int1782_t is
  variable rv : int1782_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1783_t_to_slv(x : uint1783_t) return std_logic_vector is
  variable rv : std_logic_vector(1782 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1783_t(x : std_logic_vector) return uint1783_t is
  variable rv : uint1783_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1783_t_to_slv(x : int1783_t) return std_logic_vector is
  variable rv : std_logic_vector(1782 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1783_t(x : std_logic_vector) return int1783_t is
  variable rv : int1783_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1784_t_to_slv(x : uint1784_t) return std_logic_vector is
  variable rv : std_logic_vector(1783 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1784_t(x : std_logic_vector) return uint1784_t is
  variable rv : uint1784_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1784_t_to_slv(x : int1784_t) return std_logic_vector is
  variable rv : std_logic_vector(1783 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1784_t(x : std_logic_vector) return int1784_t is
  variable rv : int1784_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1785_t_to_slv(x : uint1785_t) return std_logic_vector is
  variable rv : std_logic_vector(1784 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1785_t(x : std_logic_vector) return uint1785_t is
  variable rv : uint1785_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1785_t_to_slv(x : int1785_t) return std_logic_vector is
  variable rv : std_logic_vector(1784 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1785_t(x : std_logic_vector) return int1785_t is
  variable rv : int1785_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1786_t_to_slv(x : uint1786_t) return std_logic_vector is
  variable rv : std_logic_vector(1785 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1786_t(x : std_logic_vector) return uint1786_t is
  variable rv : uint1786_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1786_t_to_slv(x : int1786_t) return std_logic_vector is
  variable rv : std_logic_vector(1785 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1786_t(x : std_logic_vector) return int1786_t is
  variable rv : int1786_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1787_t_to_slv(x : uint1787_t) return std_logic_vector is
  variable rv : std_logic_vector(1786 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1787_t(x : std_logic_vector) return uint1787_t is
  variable rv : uint1787_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1787_t_to_slv(x : int1787_t) return std_logic_vector is
  variable rv : std_logic_vector(1786 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1787_t(x : std_logic_vector) return int1787_t is
  variable rv : int1787_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1788_t_to_slv(x : uint1788_t) return std_logic_vector is
  variable rv : std_logic_vector(1787 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1788_t(x : std_logic_vector) return uint1788_t is
  variable rv : uint1788_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1788_t_to_slv(x : int1788_t) return std_logic_vector is
  variable rv : std_logic_vector(1787 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1788_t(x : std_logic_vector) return int1788_t is
  variable rv : int1788_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1789_t_to_slv(x : uint1789_t) return std_logic_vector is
  variable rv : std_logic_vector(1788 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1789_t(x : std_logic_vector) return uint1789_t is
  variable rv : uint1789_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1789_t_to_slv(x : int1789_t) return std_logic_vector is
  variable rv : std_logic_vector(1788 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1789_t(x : std_logic_vector) return int1789_t is
  variable rv : int1789_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1790_t_to_slv(x : uint1790_t) return std_logic_vector is
  variable rv : std_logic_vector(1789 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1790_t(x : std_logic_vector) return uint1790_t is
  variable rv : uint1790_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1790_t_to_slv(x : int1790_t) return std_logic_vector is
  variable rv : std_logic_vector(1789 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1790_t(x : std_logic_vector) return int1790_t is
  variable rv : int1790_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1791_t_to_slv(x : uint1791_t) return std_logic_vector is
  variable rv : std_logic_vector(1790 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1791_t(x : std_logic_vector) return uint1791_t is
  variable rv : uint1791_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1791_t_to_slv(x : int1791_t) return std_logic_vector is
  variable rv : std_logic_vector(1790 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1791_t(x : std_logic_vector) return int1791_t is
  variable rv : int1791_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1792_t_to_slv(x : uint1792_t) return std_logic_vector is
  variable rv : std_logic_vector(1791 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1792_t(x : std_logic_vector) return uint1792_t is
  variable rv : uint1792_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1792_t_to_slv(x : int1792_t) return std_logic_vector is
  variable rv : std_logic_vector(1791 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1792_t(x : std_logic_vector) return int1792_t is
  variable rv : int1792_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1793_t_to_slv(x : uint1793_t) return std_logic_vector is
  variable rv : std_logic_vector(1792 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1793_t(x : std_logic_vector) return uint1793_t is
  variable rv : uint1793_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1793_t_to_slv(x : int1793_t) return std_logic_vector is
  variable rv : std_logic_vector(1792 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1793_t(x : std_logic_vector) return int1793_t is
  variable rv : int1793_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1794_t_to_slv(x : uint1794_t) return std_logic_vector is
  variable rv : std_logic_vector(1793 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1794_t(x : std_logic_vector) return uint1794_t is
  variable rv : uint1794_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1794_t_to_slv(x : int1794_t) return std_logic_vector is
  variable rv : std_logic_vector(1793 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1794_t(x : std_logic_vector) return int1794_t is
  variable rv : int1794_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1795_t_to_slv(x : uint1795_t) return std_logic_vector is
  variable rv : std_logic_vector(1794 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1795_t(x : std_logic_vector) return uint1795_t is
  variable rv : uint1795_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1795_t_to_slv(x : int1795_t) return std_logic_vector is
  variable rv : std_logic_vector(1794 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1795_t(x : std_logic_vector) return int1795_t is
  variable rv : int1795_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1796_t_to_slv(x : uint1796_t) return std_logic_vector is
  variable rv : std_logic_vector(1795 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1796_t(x : std_logic_vector) return uint1796_t is
  variable rv : uint1796_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1796_t_to_slv(x : int1796_t) return std_logic_vector is
  variable rv : std_logic_vector(1795 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1796_t(x : std_logic_vector) return int1796_t is
  variable rv : int1796_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1797_t_to_slv(x : uint1797_t) return std_logic_vector is
  variable rv : std_logic_vector(1796 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1797_t(x : std_logic_vector) return uint1797_t is
  variable rv : uint1797_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1797_t_to_slv(x : int1797_t) return std_logic_vector is
  variable rv : std_logic_vector(1796 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1797_t(x : std_logic_vector) return int1797_t is
  variable rv : int1797_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1798_t_to_slv(x : uint1798_t) return std_logic_vector is
  variable rv : std_logic_vector(1797 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1798_t(x : std_logic_vector) return uint1798_t is
  variable rv : uint1798_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1798_t_to_slv(x : int1798_t) return std_logic_vector is
  variable rv : std_logic_vector(1797 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1798_t(x : std_logic_vector) return int1798_t is
  variable rv : int1798_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1799_t_to_slv(x : uint1799_t) return std_logic_vector is
  variable rv : std_logic_vector(1798 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1799_t(x : std_logic_vector) return uint1799_t is
  variable rv : uint1799_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1799_t_to_slv(x : int1799_t) return std_logic_vector is
  variable rv : std_logic_vector(1798 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1799_t(x : std_logic_vector) return int1799_t is
  variable rv : int1799_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1800_t_to_slv(x : uint1800_t) return std_logic_vector is
  variable rv : std_logic_vector(1799 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1800_t(x : std_logic_vector) return uint1800_t is
  variable rv : uint1800_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1800_t_to_slv(x : int1800_t) return std_logic_vector is
  variable rv : std_logic_vector(1799 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1800_t(x : std_logic_vector) return int1800_t is
  variable rv : int1800_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1801_t_to_slv(x : uint1801_t) return std_logic_vector is
  variable rv : std_logic_vector(1800 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1801_t(x : std_logic_vector) return uint1801_t is
  variable rv : uint1801_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1801_t_to_slv(x : int1801_t) return std_logic_vector is
  variable rv : std_logic_vector(1800 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1801_t(x : std_logic_vector) return int1801_t is
  variable rv : int1801_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1802_t_to_slv(x : uint1802_t) return std_logic_vector is
  variable rv : std_logic_vector(1801 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1802_t(x : std_logic_vector) return uint1802_t is
  variable rv : uint1802_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1802_t_to_slv(x : int1802_t) return std_logic_vector is
  variable rv : std_logic_vector(1801 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1802_t(x : std_logic_vector) return int1802_t is
  variable rv : int1802_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1803_t_to_slv(x : uint1803_t) return std_logic_vector is
  variable rv : std_logic_vector(1802 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1803_t(x : std_logic_vector) return uint1803_t is
  variable rv : uint1803_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1803_t_to_slv(x : int1803_t) return std_logic_vector is
  variable rv : std_logic_vector(1802 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1803_t(x : std_logic_vector) return int1803_t is
  variable rv : int1803_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1804_t_to_slv(x : uint1804_t) return std_logic_vector is
  variable rv : std_logic_vector(1803 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1804_t(x : std_logic_vector) return uint1804_t is
  variable rv : uint1804_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1804_t_to_slv(x : int1804_t) return std_logic_vector is
  variable rv : std_logic_vector(1803 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1804_t(x : std_logic_vector) return int1804_t is
  variable rv : int1804_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1805_t_to_slv(x : uint1805_t) return std_logic_vector is
  variable rv : std_logic_vector(1804 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1805_t(x : std_logic_vector) return uint1805_t is
  variable rv : uint1805_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1805_t_to_slv(x : int1805_t) return std_logic_vector is
  variable rv : std_logic_vector(1804 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1805_t(x : std_logic_vector) return int1805_t is
  variable rv : int1805_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1806_t_to_slv(x : uint1806_t) return std_logic_vector is
  variable rv : std_logic_vector(1805 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1806_t(x : std_logic_vector) return uint1806_t is
  variable rv : uint1806_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1806_t_to_slv(x : int1806_t) return std_logic_vector is
  variable rv : std_logic_vector(1805 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1806_t(x : std_logic_vector) return int1806_t is
  variable rv : int1806_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1807_t_to_slv(x : uint1807_t) return std_logic_vector is
  variable rv : std_logic_vector(1806 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1807_t(x : std_logic_vector) return uint1807_t is
  variable rv : uint1807_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1807_t_to_slv(x : int1807_t) return std_logic_vector is
  variable rv : std_logic_vector(1806 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1807_t(x : std_logic_vector) return int1807_t is
  variable rv : int1807_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1808_t_to_slv(x : uint1808_t) return std_logic_vector is
  variable rv : std_logic_vector(1807 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1808_t(x : std_logic_vector) return uint1808_t is
  variable rv : uint1808_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1808_t_to_slv(x : int1808_t) return std_logic_vector is
  variable rv : std_logic_vector(1807 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1808_t(x : std_logic_vector) return int1808_t is
  variable rv : int1808_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1809_t_to_slv(x : uint1809_t) return std_logic_vector is
  variable rv : std_logic_vector(1808 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1809_t(x : std_logic_vector) return uint1809_t is
  variable rv : uint1809_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1809_t_to_slv(x : int1809_t) return std_logic_vector is
  variable rv : std_logic_vector(1808 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1809_t(x : std_logic_vector) return int1809_t is
  variable rv : int1809_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1810_t_to_slv(x : uint1810_t) return std_logic_vector is
  variable rv : std_logic_vector(1809 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1810_t(x : std_logic_vector) return uint1810_t is
  variable rv : uint1810_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1810_t_to_slv(x : int1810_t) return std_logic_vector is
  variable rv : std_logic_vector(1809 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1810_t(x : std_logic_vector) return int1810_t is
  variable rv : int1810_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1811_t_to_slv(x : uint1811_t) return std_logic_vector is
  variable rv : std_logic_vector(1810 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1811_t(x : std_logic_vector) return uint1811_t is
  variable rv : uint1811_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1811_t_to_slv(x : int1811_t) return std_logic_vector is
  variable rv : std_logic_vector(1810 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1811_t(x : std_logic_vector) return int1811_t is
  variable rv : int1811_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1812_t_to_slv(x : uint1812_t) return std_logic_vector is
  variable rv : std_logic_vector(1811 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1812_t(x : std_logic_vector) return uint1812_t is
  variable rv : uint1812_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1812_t_to_slv(x : int1812_t) return std_logic_vector is
  variable rv : std_logic_vector(1811 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1812_t(x : std_logic_vector) return int1812_t is
  variable rv : int1812_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1813_t_to_slv(x : uint1813_t) return std_logic_vector is
  variable rv : std_logic_vector(1812 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1813_t(x : std_logic_vector) return uint1813_t is
  variable rv : uint1813_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1813_t_to_slv(x : int1813_t) return std_logic_vector is
  variable rv : std_logic_vector(1812 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1813_t(x : std_logic_vector) return int1813_t is
  variable rv : int1813_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1814_t_to_slv(x : uint1814_t) return std_logic_vector is
  variable rv : std_logic_vector(1813 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1814_t(x : std_logic_vector) return uint1814_t is
  variable rv : uint1814_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1814_t_to_slv(x : int1814_t) return std_logic_vector is
  variable rv : std_logic_vector(1813 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1814_t(x : std_logic_vector) return int1814_t is
  variable rv : int1814_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1815_t_to_slv(x : uint1815_t) return std_logic_vector is
  variable rv : std_logic_vector(1814 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1815_t(x : std_logic_vector) return uint1815_t is
  variable rv : uint1815_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1815_t_to_slv(x : int1815_t) return std_logic_vector is
  variable rv : std_logic_vector(1814 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1815_t(x : std_logic_vector) return int1815_t is
  variable rv : int1815_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1816_t_to_slv(x : uint1816_t) return std_logic_vector is
  variable rv : std_logic_vector(1815 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1816_t(x : std_logic_vector) return uint1816_t is
  variable rv : uint1816_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1816_t_to_slv(x : int1816_t) return std_logic_vector is
  variable rv : std_logic_vector(1815 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1816_t(x : std_logic_vector) return int1816_t is
  variable rv : int1816_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1817_t_to_slv(x : uint1817_t) return std_logic_vector is
  variable rv : std_logic_vector(1816 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1817_t(x : std_logic_vector) return uint1817_t is
  variable rv : uint1817_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1817_t_to_slv(x : int1817_t) return std_logic_vector is
  variable rv : std_logic_vector(1816 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1817_t(x : std_logic_vector) return int1817_t is
  variable rv : int1817_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1818_t_to_slv(x : uint1818_t) return std_logic_vector is
  variable rv : std_logic_vector(1817 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1818_t(x : std_logic_vector) return uint1818_t is
  variable rv : uint1818_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1818_t_to_slv(x : int1818_t) return std_logic_vector is
  variable rv : std_logic_vector(1817 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1818_t(x : std_logic_vector) return int1818_t is
  variable rv : int1818_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1819_t_to_slv(x : uint1819_t) return std_logic_vector is
  variable rv : std_logic_vector(1818 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1819_t(x : std_logic_vector) return uint1819_t is
  variable rv : uint1819_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1819_t_to_slv(x : int1819_t) return std_logic_vector is
  variable rv : std_logic_vector(1818 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1819_t(x : std_logic_vector) return int1819_t is
  variable rv : int1819_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1820_t_to_slv(x : uint1820_t) return std_logic_vector is
  variable rv : std_logic_vector(1819 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1820_t(x : std_logic_vector) return uint1820_t is
  variable rv : uint1820_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1820_t_to_slv(x : int1820_t) return std_logic_vector is
  variable rv : std_logic_vector(1819 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1820_t(x : std_logic_vector) return int1820_t is
  variable rv : int1820_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1821_t_to_slv(x : uint1821_t) return std_logic_vector is
  variable rv : std_logic_vector(1820 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1821_t(x : std_logic_vector) return uint1821_t is
  variable rv : uint1821_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1821_t_to_slv(x : int1821_t) return std_logic_vector is
  variable rv : std_logic_vector(1820 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1821_t(x : std_logic_vector) return int1821_t is
  variable rv : int1821_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1822_t_to_slv(x : uint1822_t) return std_logic_vector is
  variable rv : std_logic_vector(1821 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1822_t(x : std_logic_vector) return uint1822_t is
  variable rv : uint1822_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1822_t_to_slv(x : int1822_t) return std_logic_vector is
  variable rv : std_logic_vector(1821 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1822_t(x : std_logic_vector) return int1822_t is
  variable rv : int1822_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1823_t_to_slv(x : uint1823_t) return std_logic_vector is
  variable rv : std_logic_vector(1822 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1823_t(x : std_logic_vector) return uint1823_t is
  variable rv : uint1823_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1823_t_to_slv(x : int1823_t) return std_logic_vector is
  variable rv : std_logic_vector(1822 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1823_t(x : std_logic_vector) return int1823_t is
  variable rv : int1823_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1824_t_to_slv(x : uint1824_t) return std_logic_vector is
  variable rv : std_logic_vector(1823 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1824_t(x : std_logic_vector) return uint1824_t is
  variable rv : uint1824_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1824_t_to_slv(x : int1824_t) return std_logic_vector is
  variable rv : std_logic_vector(1823 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1824_t(x : std_logic_vector) return int1824_t is
  variable rv : int1824_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1825_t_to_slv(x : uint1825_t) return std_logic_vector is
  variable rv : std_logic_vector(1824 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1825_t(x : std_logic_vector) return uint1825_t is
  variable rv : uint1825_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1825_t_to_slv(x : int1825_t) return std_logic_vector is
  variable rv : std_logic_vector(1824 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1825_t(x : std_logic_vector) return int1825_t is
  variable rv : int1825_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1826_t_to_slv(x : uint1826_t) return std_logic_vector is
  variable rv : std_logic_vector(1825 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1826_t(x : std_logic_vector) return uint1826_t is
  variable rv : uint1826_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1826_t_to_slv(x : int1826_t) return std_logic_vector is
  variable rv : std_logic_vector(1825 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1826_t(x : std_logic_vector) return int1826_t is
  variable rv : int1826_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1827_t_to_slv(x : uint1827_t) return std_logic_vector is
  variable rv : std_logic_vector(1826 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1827_t(x : std_logic_vector) return uint1827_t is
  variable rv : uint1827_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1827_t_to_slv(x : int1827_t) return std_logic_vector is
  variable rv : std_logic_vector(1826 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1827_t(x : std_logic_vector) return int1827_t is
  variable rv : int1827_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1828_t_to_slv(x : uint1828_t) return std_logic_vector is
  variable rv : std_logic_vector(1827 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1828_t(x : std_logic_vector) return uint1828_t is
  variable rv : uint1828_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1828_t_to_slv(x : int1828_t) return std_logic_vector is
  variable rv : std_logic_vector(1827 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1828_t(x : std_logic_vector) return int1828_t is
  variable rv : int1828_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1829_t_to_slv(x : uint1829_t) return std_logic_vector is
  variable rv : std_logic_vector(1828 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1829_t(x : std_logic_vector) return uint1829_t is
  variable rv : uint1829_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1829_t_to_slv(x : int1829_t) return std_logic_vector is
  variable rv : std_logic_vector(1828 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1829_t(x : std_logic_vector) return int1829_t is
  variable rv : int1829_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1830_t_to_slv(x : uint1830_t) return std_logic_vector is
  variable rv : std_logic_vector(1829 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1830_t(x : std_logic_vector) return uint1830_t is
  variable rv : uint1830_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1830_t_to_slv(x : int1830_t) return std_logic_vector is
  variable rv : std_logic_vector(1829 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1830_t(x : std_logic_vector) return int1830_t is
  variable rv : int1830_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1831_t_to_slv(x : uint1831_t) return std_logic_vector is
  variable rv : std_logic_vector(1830 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1831_t(x : std_logic_vector) return uint1831_t is
  variable rv : uint1831_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1831_t_to_slv(x : int1831_t) return std_logic_vector is
  variable rv : std_logic_vector(1830 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1831_t(x : std_logic_vector) return int1831_t is
  variable rv : int1831_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1832_t_to_slv(x : uint1832_t) return std_logic_vector is
  variable rv : std_logic_vector(1831 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1832_t(x : std_logic_vector) return uint1832_t is
  variable rv : uint1832_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1832_t_to_slv(x : int1832_t) return std_logic_vector is
  variable rv : std_logic_vector(1831 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1832_t(x : std_logic_vector) return int1832_t is
  variable rv : int1832_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1833_t_to_slv(x : uint1833_t) return std_logic_vector is
  variable rv : std_logic_vector(1832 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1833_t(x : std_logic_vector) return uint1833_t is
  variable rv : uint1833_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1833_t_to_slv(x : int1833_t) return std_logic_vector is
  variable rv : std_logic_vector(1832 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1833_t(x : std_logic_vector) return int1833_t is
  variable rv : int1833_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1834_t_to_slv(x : uint1834_t) return std_logic_vector is
  variable rv : std_logic_vector(1833 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1834_t(x : std_logic_vector) return uint1834_t is
  variable rv : uint1834_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1834_t_to_slv(x : int1834_t) return std_logic_vector is
  variable rv : std_logic_vector(1833 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1834_t(x : std_logic_vector) return int1834_t is
  variable rv : int1834_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1835_t_to_slv(x : uint1835_t) return std_logic_vector is
  variable rv : std_logic_vector(1834 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1835_t(x : std_logic_vector) return uint1835_t is
  variable rv : uint1835_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1835_t_to_slv(x : int1835_t) return std_logic_vector is
  variable rv : std_logic_vector(1834 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1835_t(x : std_logic_vector) return int1835_t is
  variable rv : int1835_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1836_t_to_slv(x : uint1836_t) return std_logic_vector is
  variable rv : std_logic_vector(1835 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1836_t(x : std_logic_vector) return uint1836_t is
  variable rv : uint1836_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1836_t_to_slv(x : int1836_t) return std_logic_vector is
  variable rv : std_logic_vector(1835 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1836_t(x : std_logic_vector) return int1836_t is
  variable rv : int1836_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1837_t_to_slv(x : uint1837_t) return std_logic_vector is
  variable rv : std_logic_vector(1836 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1837_t(x : std_logic_vector) return uint1837_t is
  variable rv : uint1837_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1837_t_to_slv(x : int1837_t) return std_logic_vector is
  variable rv : std_logic_vector(1836 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1837_t(x : std_logic_vector) return int1837_t is
  variable rv : int1837_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1838_t_to_slv(x : uint1838_t) return std_logic_vector is
  variable rv : std_logic_vector(1837 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1838_t(x : std_logic_vector) return uint1838_t is
  variable rv : uint1838_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1838_t_to_slv(x : int1838_t) return std_logic_vector is
  variable rv : std_logic_vector(1837 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1838_t(x : std_logic_vector) return int1838_t is
  variable rv : int1838_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1839_t_to_slv(x : uint1839_t) return std_logic_vector is
  variable rv : std_logic_vector(1838 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1839_t(x : std_logic_vector) return uint1839_t is
  variable rv : uint1839_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1839_t_to_slv(x : int1839_t) return std_logic_vector is
  variable rv : std_logic_vector(1838 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1839_t(x : std_logic_vector) return int1839_t is
  variable rv : int1839_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1840_t_to_slv(x : uint1840_t) return std_logic_vector is
  variable rv : std_logic_vector(1839 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1840_t(x : std_logic_vector) return uint1840_t is
  variable rv : uint1840_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1840_t_to_slv(x : int1840_t) return std_logic_vector is
  variable rv : std_logic_vector(1839 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1840_t(x : std_logic_vector) return int1840_t is
  variable rv : int1840_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1841_t_to_slv(x : uint1841_t) return std_logic_vector is
  variable rv : std_logic_vector(1840 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1841_t(x : std_logic_vector) return uint1841_t is
  variable rv : uint1841_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1841_t_to_slv(x : int1841_t) return std_logic_vector is
  variable rv : std_logic_vector(1840 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1841_t(x : std_logic_vector) return int1841_t is
  variable rv : int1841_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1842_t_to_slv(x : uint1842_t) return std_logic_vector is
  variable rv : std_logic_vector(1841 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1842_t(x : std_logic_vector) return uint1842_t is
  variable rv : uint1842_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1842_t_to_slv(x : int1842_t) return std_logic_vector is
  variable rv : std_logic_vector(1841 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1842_t(x : std_logic_vector) return int1842_t is
  variable rv : int1842_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1843_t_to_slv(x : uint1843_t) return std_logic_vector is
  variable rv : std_logic_vector(1842 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1843_t(x : std_logic_vector) return uint1843_t is
  variable rv : uint1843_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1843_t_to_slv(x : int1843_t) return std_logic_vector is
  variable rv : std_logic_vector(1842 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1843_t(x : std_logic_vector) return int1843_t is
  variable rv : int1843_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1844_t_to_slv(x : uint1844_t) return std_logic_vector is
  variable rv : std_logic_vector(1843 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1844_t(x : std_logic_vector) return uint1844_t is
  variable rv : uint1844_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1844_t_to_slv(x : int1844_t) return std_logic_vector is
  variable rv : std_logic_vector(1843 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1844_t(x : std_logic_vector) return int1844_t is
  variable rv : int1844_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1845_t_to_slv(x : uint1845_t) return std_logic_vector is
  variable rv : std_logic_vector(1844 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1845_t(x : std_logic_vector) return uint1845_t is
  variable rv : uint1845_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1845_t_to_slv(x : int1845_t) return std_logic_vector is
  variable rv : std_logic_vector(1844 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1845_t(x : std_logic_vector) return int1845_t is
  variable rv : int1845_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1846_t_to_slv(x : uint1846_t) return std_logic_vector is
  variable rv : std_logic_vector(1845 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1846_t(x : std_logic_vector) return uint1846_t is
  variable rv : uint1846_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1846_t_to_slv(x : int1846_t) return std_logic_vector is
  variable rv : std_logic_vector(1845 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1846_t(x : std_logic_vector) return int1846_t is
  variable rv : int1846_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1847_t_to_slv(x : uint1847_t) return std_logic_vector is
  variable rv : std_logic_vector(1846 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1847_t(x : std_logic_vector) return uint1847_t is
  variable rv : uint1847_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1847_t_to_slv(x : int1847_t) return std_logic_vector is
  variable rv : std_logic_vector(1846 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1847_t(x : std_logic_vector) return int1847_t is
  variable rv : int1847_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1848_t_to_slv(x : uint1848_t) return std_logic_vector is
  variable rv : std_logic_vector(1847 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1848_t(x : std_logic_vector) return uint1848_t is
  variable rv : uint1848_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1848_t_to_slv(x : int1848_t) return std_logic_vector is
  variable rv : std_logic_vector(1847 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1848_t(x : std_logic_vector) return int1848_t is
  variable rv : int1848_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1849_t_to_slv(x : uint1849_t) return std_logic_vector is
  variable rv : std_logic_vector(1848 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1849_t(x : std_logic_vector) return uint1849_t is
  variable rv : uint1849_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1849_t_to_slv(x : int1849_t) return std_logic_vector is
  variable rv : std_logic_vector(1848 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1849_t(x : std_logic_vector) return int1849_t is
  variable rv : int1849_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1850_t_to_slv(x : uint1850_t) return std_logic_vector is
  variable rv : std_logic_vector(1849 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1850_t(x : std_logic_vector) return uint1850_t is
  variable rv : uint1850_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1850_t_to_slv(x : int1850_t) return std_logic_vector is
  variable rv : std_logic_vector(1849 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1850_t(x : std_logic_vector) return int1850_t is
  variable rv : int1850_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1851_t_to_slv(x : uint1851_t) return std_logic_vector is
  variable rv : std_logic_vector(1850 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1851_t(x : std_logic_vector) return uint1851_t is
  variable rv : uint1851_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1851_t_to_slv(x : int1851_t) return std_logic_vector is
  variable rv : std_logic_vector(1850 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1851_t(x : std_logic_vector) return int1851_t is
  variable rv : int1851_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1852_t_to_slv(x : uint1852_t) return std_logic_vector is
  variable rv : std_logic_vector(1851 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1852_t(x : std_logic_vector) return uint1852_t is
  variable rv : uint1852_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1852_t_to_slv(x : int1852_t) return std_logic_vector is
  variable rv : std_logic_vector(1851 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1852_t(x : std_logic_vector) return int1852_t is
  variable rv : int1852_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1853_t_to_slv(x : uint1853_t) return std_logic_vector is
  variable rv : std_logic_vector(1852 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1853_t(x : std_logic_vector) return uint1853_t is
  variable rv : uint1853_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1853_t_to_slv(x : int1853_t) return std_logic_vector is
  variable rv : std_logic_vector(1852 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1853_t(x : std_logic_vector) return int1853_t is
  variable rv : int1853_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1854_t_to_slv(x : uint1854_t) return std_logic_vector is
  variable rv : std_logic_vector(1853 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1854_t(x : std_logic_vector) return uint1854_t is
  variable rv : uint1854_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1854_t_to_slv(x : int1854_t) return std_logic_vector is
  variable rv : std_logic_vector(1853 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1854_t(x : std_logic_vector) return int1854_t is
  variable rv : int1854_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1855_t_to_slv(x : uint1855_t) return std_logic_vector is
  variable rv : std_logic_vector(1854 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1855_t(x : std_logic_vector) return uint1855_t is
  variable rv : uint1855_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1855_t_to_slv(x : int1855_t) return std_logic_vector is
  variable rv : std_logic_vector(1854 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1855_t(x : std_logic_vector) return int1855_t is
  variable rv : int1855_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1856_t_to_slv(x : uint1856_t) return std_logic_vector is
  variable rv : std_logic_vector(1855 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1856_t(x : std_logic_vector) return uint1856_t is
  variable rv : uint1856_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1856_t_to_slv(x : int1856_t) return std_logic_vector is
  variable rv : std_logic_vector(1855 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1856_t(x : std_logic_vector) return int1856_t is
  variable rv : int1856_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1857_t_to_slv(x : uint1857_t) return std_logic_vector is
  variable rv : std_logic_vector(1856 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1857_t(x : std_logic_vector) return uint1857_t is
  variable rv : uint1857_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1857_t_to_slv(x : int1857_t) return std_logic_vector is
  variable rv : std_logic_vector(1856 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1857_t(x : std_logic_vector) return int1857_t is
  variable rv : int1857_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1858_t_to_slv(x : uint1858_t) return std_logic_vector is
  variable rv : std_logic_vector(1857 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1858_t(x : std_logic_vector) return uint1858_t is
  variable rv : uint1858_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1858_t_to_slv(x : int1858_t) return std_logic_vector is
  variable rv : std_logic_vector(1857 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1858_t(x : std_logic_vector) return int1858_t is
  variable rv : int1858_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1859_t_to_slv(x : uint1859_t) return std_logic_vector is
  variable rv : std_logic_vector(1858 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1859_t(x : std_logic_vector) return uint1859_t is
  variable rv : uint1859_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1859_t_to_slv(x : int1859_t) return std_logic_vector is
  variable rv : std_logic_vector(1858 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1859_t(x : std_logic_vector) return int1859_t is
  variable rv : int1859_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1860_t_to_slv(x : uint1860_t) return std_logic_vector is
  variable rv : std_logic_vector(1859 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1860_t(x : std_logic_vector) return uint1860_t is
  variable rv : uint1860_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1860_t_to_slv(x : int1860_t) return std_logic_vector is
  variable rv : std_logic_vector(1859 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1860_t(x : std_logic_vector) return int1860_t is
  variable rv : int1860_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1861_t_to_slv(x : uint1861_t) return std_logic_vector is
  variable rv : std_logic_vector(1860 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1861_t(x : std_logic_vector) return uint1861_t is
  variable rv : uint1861_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1861_t_to_slv(x : int1861_t) return std_logic_vector is
  variable rv : std_logic_vector(1860 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1861_t(x : std_logic_vector) return int1861_t is
  variable rv : int1861_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1862_t_to_slv(x : uint1862_t) return std_logic_vector is
  variable rv : std_logic_vector(1861 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1862_t(x : std_logic_vector) return uint1862_t is
  variable rv : uint1862_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1862_t_to_slv(x : int1862_t) return std_logic_vector is
  variable rv : std_logic_vector(1861 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1862_t(x : std_logic_vector) return int1862_t is
  variable rv : int1862_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1863_t_to_slv(x : uint1863_t) return std_logic_vector is
  variable rv : std_logic_vector(1862 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1863_t(x : std_logic_vector) return uint1863_t is
  variable rv : uint1863_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1863_t_to_slv(x : int1863_t) return std_logic_vector is
  variable rv : std_logic_vector(1862 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1863_t(x : std_logic_vector) return int1863_t is
  variable rv : int1863_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1864_t_to_slv(x : uint1864_t) return std_logic_vector is
  variable rv : std_logic_vector(1863 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1864_t(x : std_logic_vector) return uint1864_t is
  variable rv : uint1864_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1864_t_to_slv(x : int1864_t) return std_logic_vector is
  variable rv : std_logic_vector(1863 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1864_t(x : std_logic_vector) return int1864_t is
  variable rv : int1864_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1865_t_to_slv(x : uint1865_t) return std_logic_vector is
  variable rv : std_logic_vector(1864 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1865_t(x : std_logic_vector) return uint1865_t is
  variable rv : uint1865_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1865_t_to_slv(x : int1865_t) return std_logic_vector is
  variable rv : std_logic_vector(1864 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1865_t(x : std_logic_vector) return int1865_t is
  variable rv : int1865_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1866_t_to_slv(x : uint1866_t) return std_logic_vector is
  variable rv : std_logic_vector(1865 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1866_t(x : std_logic_vector) return uint1866_t is
  variable rv : uint1866_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1866_t_to_slv(x : int1866_t) return std_logic_vector is
  variable rv : std_logic_vector(1865 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1866_t(x : std_logic_vector) return int1866_t is
  variable rv : int1866_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1867_t_to_slv(x : uint1867_t) return std_logic_vector is
  variable rv : std_logic_vector(1866 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1867_t(x : std_logic_vector) return uint1867_t is
  variable rv : uint1867_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1867_t_to_slv(x : int1867_t) return std_logic_vector is
  variable rv : std_logic_vector(1866 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1867_t(x : std_logic_vector) return int1867_t is
  variable rv : int1867_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1868_t_to_slv(x : uint1868_t) return std_logic_vector is
  variable rv : std_logic_vector(1867 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1868_t(x : std_logic_vector) return uint1868_t is
  variable rv : uint1868_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1868_t_to_slv(x : int1868_t) return std_logic_vector is
  variable rv : std_logic_vector(1867 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1868_t(x : std_logic_vector) return int1868_t is
  variable rv : int1868_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1869_t_to_slv(x : uint1869_t) return std_logic_vector is
  variable rv : std_logic_vector(1868 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1869_t(x : std_logic_vector) return uint1869_t is
  variable rv : uint1869_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1869_t_to_slv(x : int1869_t) return std_logic_vector is
  variable rv : std_logic_vector(1868 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1869_t(x : std_logic_vector) return int1869_t is
  variable rv : int1869_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1870_t_to_slv(x : uint1870_t) return std_logic_vector is
  variable rv : std_logic_vector(1869 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1870_t(x : std_logic_vector) return uint1870_t is
  variable rv : uint1870_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1870_t_to_slv(x : int1870_t) return std_logic_vector is
  variable rv : std_logic_vector(1869 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1870_t(x : std_logic_vector) return int1870_t is
  variable rv : int1870_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1871_t_to_slv(x : uint1871_t) return std_logic_vector is
  variable rv : std_logic_vector(1870 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1871_t(x : std_logic_vector) return uint1871_t is
  variable rv : uint1871_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1871_t_to_slv(x : int1871_t) return std_logic_vector is
  variable rv : std_logic_vector(1870 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1871_t(x : std_logic_vector) return int1871_t is
  variable rv : int1871_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1872_t_to_slv(x : uint1872_t) return std_logic_vector is
  variable rv : std_logic_vector(1871 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1872_t(x : std_logic_vector) return uint1872_t is
  variable rv : uint1872_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1872_t_to_slv(x : int1872_t) return std_logic_vector is
  variable rv : std_logic_vector(1871 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1872_t(x : std_logic_vector) return int1872_t is
  variable rv : int1872_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1873_t_to_slv(x : uint1873_t) return std_logic_vector is
  variable rv : std_logic_vector(1872 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1873_t(x : std_logic_vector) return uint1873_t is
  variable rv : uint1873_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1873_t_to_slv(x : int1873_t) return std_logic_vector is
  variable rv : std_logic_vector(1872 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1873_t(x : std_logic_vector) return int1873_t is
  variable rv : int1873_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1874_t_to_slv(x : uint1874_t) return std_logic_vector is
  variable rv : std_logic_vector(1873 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1874_t(x : std_logic_vector) return uint1874_t is
  variable rv : uint1874_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1874_t_to_slv(x : int1874_t) return std_logic_vector is
  variable rv : std_logic_vector(1873 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1874_t(x : std_logic_vector) return int1874_t is
  variable rv : int1874_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1875_t_to_slv(x : uint1875_t) return std_logic_vector is
  variable rv : std_logic_vector(1874 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1875_t(x : std_logic_vector) return uint1875_t is
  variable rv : uint1875_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1875_t_to_slv(x : int1875_t) return std_logic_vector is
  variable rv : std_logic_vector(1874 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1875_t(x : std_logic_vector) return int1875_t is
  variable rv : int1875_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1876_t_to_slv(x : uint1876_t) return std_logic_vector is
  variable rv : std_logic_vector(1875 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1876_t(x : std_logic_vector) return uint1876_t is
  variable rv : uint1876_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1876_t_to_slv(x : int1876_t) return std_logic_vector is
  variable rv : std_logic_vector(1875 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1876_t(x : std_logic_vector) return int1876_t is
  variable rv : int1876_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1877_t_to_slv(x : uint1877_t) return std_logic_vector is
  variable rv : std_logic_vector(1876 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1877_t(x : std_logic_vector) return uint1877_t is
  variable rv : uint1877_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1877_t_to_slv(x : int1877_t) return std_logic_vector is
  variable rv : std_logic_vector(1876 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1877_t(x : std_logic_vector) return int1877_t is
  variable rv : int1877_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1878_t_to_slv(x : uint1878_t) return std_logic_vector is
  variable rv : std_logic_vector(1877 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1878_t(x : std_logic_vector) return uint1878_t is
  variable rv : uint1878_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1878_t_to_slv(x : int1878_t) return std_logic_vector is
  variable rv : std_logic_vector(1877 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1878_t(x : std_logic_vector) return int1878_t is
  variable rv : int1878_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1879_t_to_slv(x : uint1879_t) return std_logic_vector is
  variable rv : std_logic_vector(1878 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1879_t(x : std_logic_vector) return uint1879_t is
  variable rv : uint1879_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1879_t_to_slv(x : int1879_t) return std_logic_vector is
  variable rv : std_logic_vector(1878 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1879_t(x : std_logic_vector) return int1879_t is
  variable rv : int1879_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1880_t_to_slv(x : uint1880_t) return std_logic_vector is
  variable rv : std_logic_vector(1879 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1880_t(x : std_logic_vector) return uint1880_t is
  variable rv : uint1880_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1880_t_to_slv(x : int1880_t) return std_logic_vector is
  variable rv : std_logic_vector(1879 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1880_t(x : std_logic_vector) return int1880_t is
  variable rv : int1880_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1881_t_to_slv(x : uint1881_t) return std_logic_vector is
  variable rv : std_logic_vector(1880 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1881_t(x : std_logic_vector) return uint1881_t is
  variable rv : uint1881_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1881_t_to_slv(x : int1881_t) return std_logic_vector is
  variable rv : std_logic_vector(1880 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1881_t(x : std_logic_vector) return int1881_t is
  variable rv : int1881_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1882_t_to_slv(x : uint1882_t) return std_logic_vector is
  variable rv : std_logic_vector(1881 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1882_t(x : std_logic_vector) return uint1882_t is
  variable rv : uint1882_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1882_t_to_slv(x : int1882_t) return std_logic_vector is
  variable rv : std_logic_vector(1881 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1882_t(x : std_logic_vector) return int1882_t is
  variable rv : int1882_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1883_t_to_slv(x : uint1883_t) return std_logic_vector is
  variable rv : std_logic_vector(1882 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1883_t(x : std_logic_vector) return uint1883_t is
  variable rv : uint1883_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1883_t_to_slv(x : int1883_t) return std_logic_vector is
  variable rv : std_logic_vector(1882 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1883_t(x : std_logic_vector) return int1883_t is
  variable rv : int1883_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1884_t_to_slv(x : uint1884_t) return std_logic_vector is
  variable rv : std_logic_vector(1883 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1884_t(x : std_logic_vector) return uint1884_t is
  variable rv : uint1884_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1884_t_to_slv(x : int1884_t) return std_logic_vector is
  variable rv : std_logic_vector(1883 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1884_t(x : std_logic_vector) return int1884_t is
  variable rv : int1884_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1885_t_to_slv(x : uint1885_t) return std_logic_vector is
  variable rv : std_logic_vector(1884 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1885_t(x : std_logic_vector) return uint1885_t is
  variable rv : uint1885_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1885_t_to_slv(x : int1885_t) return std_logic_vector is
  variable rv : std_logic_vector(1884 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1885_t(x : std_logic_vector) return int1885_t is
  variable rv : int1885_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1886_t_to_slv(x : uint1886_t) return std_logic_vector is
  variable rv : std_logic_vector(1885 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1886_t(x : std_logic_vector) return uint1886_t is
  variable rv : uint1886_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1886_t_to_slv(x : int1886_t) return std_logic_vector is
  variable rv : std_logic_vector(1885 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1886_t(x : std_logic_vector) return int1886_t is
  variable rv : int1886_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1887_t_to_slv(x : uint1887_t) return std_logic_vector is
  variable rv : std_logic_vector(1886 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1887_t(x : std_logic_vector) return uint1887_t is
  variable rv : uint1887_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1887_t_to_slv(x : int1887_t) return std_logic_vector is
  variable rv : std_logic_vector(1886 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1887_t(x : std_logic_vector) return int1887_t is
  variable rv : int1887_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1888_t_to_slv(x : uint1888_t) return std_logic_vector is
  variable rv : std_logic_vector(1887 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1888_t(x : std_logic_vector) return uint1888_t is
  variable rv : uint1888_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1888_t_to_slv(x : int1888_t) return std_logic_vector is
  variable rv : std_logic_vector(1887 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1888_t(x : std_logic_vector) return int1888_t is
  variable rv : int1888_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1889_t_to_slv(x : uint1889_t) return std_logic_vector is
  variable rv : std_logic_vector(1888 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1889_t(x : std_logic_vector) return uint1889_t is
  variable rv : uint1889_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1889_t_to_slv(x : int1889_t) return std_logic_vector is
  variable rv : std_logic_vector(1888 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1889_t(x : std_logic_vector) return int1889_t is
  variable rv : int1889_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1890_t_to_slv(x : uint1890_t) return std_logic_vector is
  variable rv : std_logic_vector(1889 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1890_t(x : std_logic_vector) return uint1890_t is
  variable rv : uint1890_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1890_t_to_slv(x : int1890_t) return std_logic_vector is
  variable rv : std_logic_vector(1889 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1890_t(x : std_logic_vector) return int1890_t is
  variable rv : int1890_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1891_t_to_slv(x : uint1891_t) return std_logic_vector is
  variable rv : std_logic_vector(1890 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1891_t(x : std_logic_vector) return uint1891_t is
  variable rv : uint1891_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1891_t_to_slv(x : int1891_t) return std_logic_vector is
  variable rv : std_logic_vector(1890 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1891_t(x : std_logic_vector) return int1891_t is
  variable rv : int1891_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1892_t_to_slv(x : uint1892_t) return std_logic_vector is
  variable rv : std_logic_vector(1891 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1892_t(x : std_logic_vector) return uint1892_t is
  variable rv : uint1892_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1892_t_to_slv(x : int1892_t) return std_logic_vector is
  variable rv : std_logic_vector(1891 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1892_t(x : std_logic_vector) return int1892_t is
  variable rv : int1892_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1893_t_to_slv(x : uint1893_t) return std_logic_vector is
  variable rv : std_logic_vector(1892 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1893_t(x : std_logic_vector) return uint1893_t is
  variable rv : uint1893_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1893_t_to_slv(x : int1893_t) return std_logic_vector is
  variable rv : std_logic_vector(1892 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1893_t(x : std_logic_vector) return int1893_t is
  variable rv : int1893_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1894_t_to_slv(x : uint1894_t) return std_logic_vector is
  variable rv : std_logic_vector(1893 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1894_t(x : std_logic_vector) return uint1894_t is
  variable rv : uint1894_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1894_t_to_slv(x : int1894_t) return std_logic_vector is
  variable rv : std_logic_vector(1893 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1894_t(x : std_logic_vector) return int1894_t is
  variable rv : int1894_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1895_t_to_slv(x : uint1895_t) return std_logic_vector is
  variable rv : std_logic_vector(1894 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1895_t(x : std_logic_vector) return uint1895_t is
  variable rv : uint1895_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1895_t_to_slv(x : int1895_t) return std_logic_vector is
  variable rv : std_logic_vector(1894 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1895_t(x : std_logic_vector) return int1895_t is
  variable rv : int1895_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1896_t_to_slv(x : uint1896_t) return std_logic_vector is
  variable rv : std_logic_vector(1895 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1896_t(x : std_logic_vector) return uint1896_t is
  variable rv : uint1896_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1896_t_to_slv(x : int1896_t) return std_logic_vector is
  variable rv : std_logic_vector(1895 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1896_t(x : std_logic_vector) return int1896_t is
  variable rv : int1896_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1897_t_to_slv(x : uint1897_t) return std_logic_vector is
  variable rv : std_logic_vector(1896 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1897_t(x : std_logic_vector) return uint1897_t is
  variable rv : uint1897_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1897_t_to_slv(x : int1897_t) return std_logic_vector is
  variable rv : std_logic_vector(1896 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1897_t(x : std_logic_vector) return int1897_t is
  variable rv : int1897_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1898_t_to_slv(x : uint1898_t) return std_logic_vector is
  variable rv : std_logic_vector(1897 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1898_t(x : std_logic_vector) return uint1898_t is
  variable rv : uint1898_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1898_t_to_slv(x : int1898_t) return std_logic_vector is
  variable rv : std_logic_vector(1897 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1898_t(x : std_logic_vector) return int1898_t is
  variable rv : int1898_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1899_t_to_slv(x : uint1899_t) return std_logic_vector is
  variable rv : std_logic_vector(1898 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1899_t(x : std_logic_vector) return uint1899_t is
  variable rv : uint1899_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1899_t_to_slv(x : int1899_t) return std_logic_vector is
  variable rv : std_logic_vector(1898 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1899_t(x : std_logic_vector) return int1899_t is
  variable rv : int1899_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1900_t_to_slv(x : uint1900_t) return std_logic_vector is
  variable rv : std_logic_vector(1899 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1900_t(x : std_logic_vector) return uint1900_t is
  variable rv : uint1900_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1900_t_to_slv(x : int1900_t) return std_logic_vector is
  variable rv : std_logic_vector(1899 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1900_t(x : std_logic_vector) return int1900_t is
  variable rv : int1900_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1901_t_to_slv(x : uint1901_t) return std_logic_vector is
  variable rv : std_logic_vector(1900 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1901_t(x : std_logic_vector) return uint1901_t is
  variable rv : uint1901_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1901_t_to_slv(x : int1901_t) return std_logic_vector is
  variable rv : std_logic_vector(1900 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1901_t(x : std_logic_vector) return int1901_t is
  variable rv : int1901_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1902_t_to_slv(x : uint1902_t) return std_logic_vector is
  variable rv : std_logic_vector(1901 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1902_t(x : std_logic_vector) return uint1902_t is
  variable rv : uint1902_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1902_t_to_slv(x : int1902_t) return std_logic_vector is
  variable rv : std_logic_vector(1901 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1902_t(x : std_logic_vector) return int1902_t is
  variable rv : int1902_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1903_t_to_slv(x : uint1903_t) return std_logic_vector is
  variable rv : std_logic_vector(1902 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1903_t(x : std_logic_vector) return uint1903_t is
  variable rv : uint1903_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1903_t_to_slv(x : int1903_t) return std_logic_vector is
  variable rv : std_logic_vector(1902 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1903_t(x : std_logic_vector) return int1903_t is
  variable rv : int1903_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1904_t_to_slv(x : uint1904_t) return std_logic_vector is
  variable rv : std_logic_vector(1903 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1904_t(x : std_logic_vector) return uint1904_t is
  variable rv : uint1904_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1904_t_to_slv(x : int1904_t) return std_logic_vector is
  variable rv : std_logic_vector(1903 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1904_t(x : std_logic_vector) return int1904_t is
  variable rv : int1904_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1905_t_to_slv(x : uint1905_t) return std_logic_vector is
  variable rv : std_logic_vector(1904 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1905_t(x : std_logic_vector) return uint1905_t is
  variable rv : uint1905_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1905_t_to_slv(x : int1905_t) return std_logic_vector is
  variable rv : std_logic_vector(1904 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1905_t(x : std_logic_vector) return int1905_t is
  variable rv : int1905_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1906_t_to_slv(x : uint1906_t) return std_logic_vector is
  variable rv : std_logic_vector(1905 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1906_t(x : std_logic_vector) return uint1906_t is
  variable rv : uint1906_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1906_t_to_slv(x : int1906_t) return std_logic_vector is
  variable rv : std_logic_vector(1905 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1906_t(x : std_logic_vector) return int1906_t is
  variable rv : int1906_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1907_t_to_slv(x : uint1907_t) return std_logic_vector is
  variable rv : std_logic_vector(1906 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1907_t(x : std_logic_vector) return uint1907_t is
  variable rv : uint1907_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1907_t_to_slv(x : int1907_t) return std_logic_vector is
  variable rv : std_logic_vector(1906 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1907_t(x : std_logic_vector) return int1907_t is
  variable rv : int1907_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1908_t_to_slv(x : uint1908_t) return std_logic_vector is
  variable rv : std_logic_vector(1907 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1908_t(x : std_logic_vector) return uint1908_t is
  variable rv : uint1908_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1908_t_to_slv(x : int1908_t) return std_logic_vector is
  variable rv : std_logic_vector(1907 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1908_t(x : std_logic_vector) return int1908_t is
  variable rv : int1908_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1909_t_to_slv(x : uint1909_t) return std_logic_vector is
  variable rv : std_logic_vector(1908 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1909_t(x : std_logic_vector) return uint1909_t is
  variable rv : uint1909_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1909_t_to_slv(x : int1909_t) return std_logic_vector is
  variable rv : std_logic_vector(1908 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1909_t(x : std_logic_vector) return int1909_t is
  variable rv : int1909_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1910_t_to_slv(x : uint1910_t) return std_logic_vector is
  variable rv : std_logic_vector(1909 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1910_t(x : std_logic_vector) return uint1910_t is
  variable rv : uint1910_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1910_t_to_slv(x : int1910_t) return std_logic_vector is
  variable rv : std_logic_vector(1909 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1910_t(x : std_logic_vector) return int1910_t is
  variable rv : int1910_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1911_t_to_slv(x : uint1911_t) return std_logic_vector is
  variable rv : std_logic_vector(1910 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1911_t(x : std_logic_vector) return uint1911_t is
  variable rv : uint1911_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1911_t_to_slv(x : int1911_t) return std_logic_vector is
  variable rv : std_logic_vector(1910 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1911_t(x : std_logic_vector) return int1911_t is
  variable rv : int1911_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1912_t_to_slv(x : uint1912_t) return std_logic_vector is
  variable rv : std_logic_vector(1911 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1912_t(x : std_logic_vector) return uint1912_t is
  variable rv : uint1912_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1912_t_to_slv(x : int1912_t) return std_logic_vector is
  variable rv : std_logic_vector(1911 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1912_t(x : std_logic_vector) return int1912_t is
  variable rv : int1912_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1913_t_to_slv(x : uint1913_t) return std_logic_vector is
  variable rv : std_logic_vector(1912 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1913_t(x : std_logic_vector) return uint1913_t is
  variable rv : uint1913_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1913_t_to_slv(x : int1913_t) return std_logic_vector is
  variable rv : std_logic_vector(1912 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1913_t(x : std_logic_vector) return int1913_t is
  variable rv : int1913_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1914_t_to_slv(x : uint1914_t) return std_logic_vector is
  variable rv : std_logic_vector(1913 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1914_t(x : std_logic_vector) return uint1914_t is
  variable rv : uint1914_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1914_t_to_slv(x : int1914_t) return std_logic_vector is
  variable rv : std_logic_vector(1913 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1914_t(x : std_logic_vector) return int1914_t is
  variable rv : int1914_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1915_t_to_slv(x : uint1915_t) return std_logic_vector is
  variable rv : std_logic_vector(1914 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1915_t(x : std_logic_vector) return uint1915_t is
  variable rv : uint1915_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1915_t_to_slv(x : int1915_t) return std_logic_vector is
  variable rv : std_logic_vector(1914 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1915_t(x : std_logic_vector) return int1915_t is
  variable rv : int1915_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1916_t_to_slv(x : uint1916_t) return std_logic_vector is
  variable rv : std_logic_vector(1915 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1916_t(x : std_logic_vector) return uint1916_t is
  variable rv : uint1916_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1916_t_to_slv(x : int1916_t) return std_logic_vector is
  variable rv : std_logic_vector(1915 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1916_t(x : std_logic_vector) return int1916_t is
  variable rv : int1916_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1917_t_to_slv(x : uint1917_t) return std_logic_vector is
  variable rv : std_logic_vector(1916 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1917_t(x : std_logic_vector) return uint1917_t is
  variable rv : uint1917_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1917_t_to_slv(x : int1917_t) return std_logic_vector is
  variable rv : std_logic_vector(1916 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1917_t(x : std_logic_vector) return int1917_t is
  variable rv : int1917_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1918_t_to_slv(x : uint1918_t) return std_logic_vector is
  variable rv : std_logic_vector(1917 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1918_t(x : std_logic_vector) return uint1918_t is
  variable rv : uint1918_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1918_t_to_slv(x : int1918_t) return std_logic_vector is
  variable rv : std_logic_vector(1917 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1918_t(x : std_logic_vector) return int1918_t is
  variable rv : int1918_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1919_t_to_slv(x : uint1919_t) return std_logic_vector is
  variable rv : std_logic_vector(1918 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1919_t(x : std_logic_vector) return uint1919_t is
  variable rv : uint1919_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1919_t_to_slv(x : int1919_t) return std_logic_vector is
  variable rv : std_logic_vector(1918 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1919_t(x : std_logic_vector) return int1919_t is
  variable rv : int1919_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1920_t_to_slv(x : uint1920_t) return std_logic_vector is
  variable rv : std_logic_vector(1919 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1920_t(x : std_logic_vector) return uint1920_t is
  variable rv : uint1920_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1920_t_to_slv(x : int1920_t) return std_logic_vector is
  variable rv : std_logic_vector(1919 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1920_t(x : std_logic_vector) return int1920_t is
  variable rv : int1920_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1921_t_to_slv(x : uint1921_t) return std_logic_vector is
  variable rv : std_logic_vector(1920 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1921_t(x : std_logic_vector) return uint1921_t is
  variable rv : uint1921_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1921_t_to_slv(x : int1921_t) return std_logic_vector is
  variable rv : std_logic_vector(1920 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1921_t(x : std_logic_vector) return int1921_t is
  variable rv : int1921_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1922_t_to_slv(x : uint1922_t) return std_logic_vector is
  variable rv : std_logic_vector(1921 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1922_t(x : std_logic_vector) return uint1922_t is
  variable rv : uint1922_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1922_t_to_slv(x : int1922_t) return std_logic_vector is
  variable rv : std_logic_vector(1921 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1922_t(x : std_logic_vector) return int1922_t is
  variable rv : int1922_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1923_t_to_slv(x : uint1923_t) return std_logic_vector is
  variable rv : std_logic_vector(1922 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1923_t(x : std_logic_vector) return uint1923_t is
  variable rv : uint1923_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1923_t_to_slv(x : int1923_t) return std_logic_vector is
  variable rv : std_logic_vector(1922 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1923_t(x : std_logic_vector) return int1923_t is
  variable rv : int1923_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1924_t_to_slv(x : uint1924_t) return std_logic_vector is
  variable rv : std_logic_vector(1923 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1924_t(x : std_logic_vector) return uint1924_t is
  variable rv : uint1924_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1924_t_to_slv(x : int1924_t) return std_logic_vector is
  variable rv : std_logic_vector(1923 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1924_t(x : std_logic_vector) return int1924_t is
  variable rv : int1924_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1925_t_to_slv(x : uint1925_t) return std_logic_vector is
  variable rv : std_logic_vector(1924 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1925_t(x : std_logic_vector) return uint1925_t is
  variable rv : uint1925_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1925_t_to_slv(x : int1925_t) return std_logic_vector is
  variable rv : std_logic_vector(1924 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1925_t(x : std_logic_vector) return int1925_t is
  variable rv : int1925_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1926_t_to_slv(x : uint1926_t) return std_logic_vector is
  variable rv : std_logic_vector(1925 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1926_t(x : std_logic_vector) return uint1926_t is
  variable rv : uint1926_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1926_t_to_slv(x : int1926_t) return std_logic_vector is
  variable rv : std_logic_vector(1925 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1926_t(x : std_logic_vector) return int1926_t is
  variable rv : int1926_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1927_t_to_slv(x : uint1927_t) return std_logic_vector is
  variable rv : std_logic_vector(1926 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1927_t(x : std_logic_vector) return uint1927_t is
  variable rv : uint1927_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1927_t_to_slv(x : int1927_t) return std_logic_vector is
  variable rv : std_logic_vector(1926 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1927_t(x : std_logic_vector) return int1927_t is
  variable rv : int1927_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1928_t_to_slv(x : uint1928_t) return std_logic_vector is
  variable rv : std_logic_vector(1927 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1928_t(x : std_logic_vector) return uint1928_t is
  variable rv : uint1928_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1928_t_to_slv(x : int1928_t) return std_logic_vector is
  variable rv : std_logic_vector(1927 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1928_t(x : std_logic_vector) return int1928_t is
  variable rv : int1928_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1929_t_to_slv(x : uint1929_t) return std_logic_vector is
  variable rv : std_logic_vector(1928 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1929_t(x : std_logic_vector) return uint1929_t is
  variable rv : uint1929_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1929_t_to_slv(x : int1929_t) return std_logic_vector is
  variable rv : std_logic_vector(1928 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1929_t(x : std_logic_vector) return int1929_t is
  variable rv : int1929_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1930_t_to_slv(x : uint1930_t) return std_logic_vector is
  variable rv : std_logic_vector(1929 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1930_t(x : std_logic_vector) return uint1930_t is
  variable rv : uint1930_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1930_t_to_slv(x : int1930_t) return std_logic_vector is
  variable rv : std_logic_vector(1929 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1930_t(x : std_logic_vector) return int1930_t is
  variable rv : int1930_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1931_t_to_slv(x : uint1931_t) return std_logic_vector is
  variable rv : std_logic_vector(1930 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1931_t(x : std_logic_vector) return uint1931_t is
  variable rv : uint1931_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1931_t_to_slv(x : int1931_t) return std_logic_vector is
  variable rv : std_logic_vector(1930 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1931_t(x : std_logic_vector) return int1931_t is
  variable rv : int1931_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1932_t_to_slv(x : uint1932_t) return std_logic_vector is
  variable rv : std_logic_vector(1931 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1932_t(x : std_logic_vector) return uint1932_t is
  variable rv : uint1932_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1932_t_to_slv(x : int1932_t) return std_logic_vector is
  variable rv : std_logic_vector(1931 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1932_t(x : std_logic_vector) return int1932_t is
  variable rv : int1932_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1933_t_to_slv(x : uint1933_t) return std_logic_vector is
  variable rv : std_logic_vector(1932 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1933_t(x : std_logic_vector) return uint1933_t is
  variable rv : uint1933_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1933_t_to_slv(x : int1933_t) return std_logic_vector is
  variable rv : std_logic_vector(1932 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1933_t(x : std_logic_vector) return int1933_t is
  variable rv : int1933_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1934_t_to_slv(x : uint1934_t) return std_logic_vector is
  variable rv : std_logic_vector(1933 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1934_t(x : std_logic_vector) return uint1934_t is
  variable rv : uint1934_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1934_t_to_slv(x : int1934_t) return std_logic_vector is
  variable rv : std_logic_vector(1933 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1934_t(x : std_logic_vector) return int1934_t is
  variable rv : int1934_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1935_t_to_slv(x : uint1935_t) return std_logic_vector is
  variable rv : std_logic_vector(1934 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1935_t(x : std_logic_vector) return uint1935_t is
  variable rv : uint1935_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1935_t_to_slv(x : int1935_t) return std_logic_vector is
  variable rv : std_logic_vector(1934 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1935_t(x : std_logic_vector) return int1935_t is
  variable rv : int1935_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1936_t_to_slv(x : uint1936_t) return std_logic_vector is
  variable rv : std_logic_vector(1935 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1936_t(x : std_logic_vector) return uint1936_t is
  variable rv : uint1936_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1936_t_to_slv(x : int1936_t) return std_logic_vector is
  variable rv : std_logic_vector(1935 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1936_t(x : std_logic_vector) return int1936_t is
  variable rv : int1936_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1937_t_to_slv(x : uint1937_t) return std_logic_vector is
  variable rv : std_logic_vector(1936 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1937_t(x : std_logic_vector) return uint1937_t is
  variable rv : uint1937_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1937_t_to_slv(x : int1937_t) return std_logic_vector is
  variable rv : std_logic_vector(1936 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1937_t(x : std_logic_vector) return int1937_t is
  variable rv : int1937_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1938_t_to_slv(x : uint1938_t) return std_logic_vector is
  variable rv : std_logic_vector(1937 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1938_t(x : std_logic_vector) return uint1938_t is
  variable rv : uint1938_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1938_t_to_slv(x : int1938_t) return std_logic_vector is
  variable rv : std_logic_vector(1937 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1938_t(x : std_logic_vector) return int1938_t is
  variable rv : int1938_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1939_t_to_slv(x : uint1939_t) return std_logic_vector is
  variable rv : std_logic_vector(1938 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1939_t(x : std_logic_vector) return uint1939_t is
  variable rv : uint1939_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1939_t_to_slv(x : int1939_t) return std_logic_vector is
  variable rv : std_logic_vector(1938 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1939_t(x : std_logic_vector) return int1939_t is
  variable rv : int1939_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1940_t_to_slv(x : uint1940_t) return std_logic_vector is
  variable rv : std_logic_vector(1939 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1940_t(x : std_logic_vector) return uint1940_t is
  variable rv : uint1940_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1940_t_to_slv(x : int1940_t) return std_logic_vector is
  variable rv : std_logic_vector(1939 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1940_t(x : std_logic_vector) return int1940_t is
  variable rv : int1940_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1941_t_to_slv(x : uint1941_t) return std_logic_vector is
  variable rv : std_logic_vector(1940 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1941_t(x : std_logic_vector) return uint1941_t is
  variable rv : uint1941_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1941_t_to_slv(x : int1941_t) return std_logic_vector is
  variable rv : std_logic_vector(1940 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1941_t(x : std_logic_vector) return int1941_t is
  variable rv : int1941_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1942_t_to_slv(x : uint1942_t) return std_logic_vector is
  variable rv : std_logic_vector(1941 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1942_t(x : std_logic_vector) return uint1942_t is
  variable rv : uint1942_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1942_t_to_slv(x : int1942_t) return std_logic_vector is
  variable rv : std_logic_vector(1941 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1942_t(x : std_logic_vector) return int1942_t is
  variable rv : int1942_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1943_t_to_slv(x : uint1943_t) return std_logic_vector is
  variable rv : std_logic_vector(1942 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1943_t(x : std_logic_vector) return uint1943_t is
  variable rv : uint1943_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1943_t_to_slv(x : int1943_t) return std_logic_vector is
  variable rv : std_logic_vector(1942 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1943_t(x : std_logic_vector) return int1943_t is
  variable rv : int1943_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1944_t_to_slv(x : uint1944_t) return std_logic_vector is
  variable rv : std_logic_vector(1943 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1944_t(x : std_logic_vector) return uint1944_t is
  variable rv : uint1944_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1944_t_to_slv(x : int1944_t) return std_logic_vector is
  variable rv : std_logic_vector(1943 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1944_t(x : std_logic_vector) return int1944_t is
  variable rv : int1944_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1945_t_to_slv(x : uint1945_t) return std_logic_vector is
  variable rv : std_logic_vector(1944 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1945_t(x : std_logic_vector) return uint1945_t is
  variable rv : uint1945_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1945_t_to_slv(x : int1945_t) return std_logic_vector is
  variable rv : std_logic_vector(1944 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1945_t(x : std_logic_vector) return int1945_t is
  variable rv : int1945_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1946_t_to_slv(x : uint1946_t) return std_logic_vector is
  variable rv : std_logic_vector(1945 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1946_t(x : std_logic_vector) return uint1946_t is
  variable rv : uint1946_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1946_t_to_slv(x : int1946_t) return std_logic_vector is
  variable rv : std_logic_vector(1945 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1946_t(x : std_logic_vector) return int1946_t is
  variable rv : int1946_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1947_t_to_slv(x : uint1947_t) return std_logic_vector is
  variable rv : std_logic_vector(1946 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1947_t(x : std_logic_vector) return uint1947_t is
  variable rv : uint1947_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1947_t_to_slv(x : int1947_t) return std_logic_vector is
  variable rv : std_logic_vector(1946 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1947_t(x : std_logic_vector) return int1947_t is
  variable rv : int1947_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1948_t_to_slv(x : uint1948_t) return std_logic_vector is
  variable rv : std_logic_vector(1947 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1948_t(x : std_logic_vector) return uint1948_t is
  variable rv : uint1948_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1948_t_to_slv(x : int1948_t) return std_logic_vector is
  variable rv : std_logic_vector(1947 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1948_t(x : std_logic_vector) return int1948_t is
  variable rv : int1948_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1949_t_to_slv(x : uint1949_t) return std_logic_vector is
  variable rv : std_logic_vector(1948 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1949_t(x : std_logic_vector) return uint1949_t is
  variable rv : uint1949_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1949_t_to_slv(x : int1949_t) return std_logic_vector is
  variable rv : std_logic_vector(1948 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1949_t(x : std_logic_vector) return int1949_t is
  variable rv : int1949_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1950_t_to_slv(x : uint1950_t) return std_logic_vector is
  variable rv : std_logic_vector(1949 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1950_t(x : std_logic_vector) return uint1950_t is
  variable rv : uint1950_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1950_t_to_slv(x : int1950_t) return std_logic_vector is
  variable rv : std_logic_vector(1949 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1950_t(x : std_logic_vector) return int1950_t is
  variable rv : int1950_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1951_t_to_slv(x : uint1951_t) return std_logic_vector is
  variable rv : std_logic_vector(1950 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1951_t(x : std_logic_vector) return uint1951_t is
  variable rv : uint1951_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1951_t_to_slv(x : int1951_t) return std_logic_vector is
  variable rv : std_logic_vector(1950 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1951_t(x : std_logic_vector) return int1951_t is
  variable rv : int1951_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1952_t_to_slv(x : uint1952_t) return std_logic_vector is
  variable rv : std_logic_vector(1951 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1952_t(x : std_logic_vector) return uint1952_t is
  variable rv : uint1952_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1952_t_to_slv(x : int1952_t) return std_logic_vector is
  variable rv : std_logic_vector(1951 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1952_t(x : std_logic_vector) return int1952_t is
  variable rv : int1952_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1953_t_to_slv(x : uint1953_t) return std_logic_vector is
  variable rv : std_logic_vector(1952 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1953_t(x : std_logic_vector) return uint1953_t is
  variable rv : uint1953_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1953_t_to_slv(x : int1953_t) return std_logic_vector is
  variable rv : std_logic_vector(1952 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1953_t(x : std_logic_vector) return int1953_t is
  variable rv : int1953_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1954_t_to_slv(x : uint1954_t) return std_logic_vector is
  variable rv : std_logic_vector(1953 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1954_t(x : std_logic_vector) return uint1954_t is
  variable rv : uint1954_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1954_t_to_slv(x : int1954_t) return std_logic_vector is
  variable rv : std_logic_vector(1953 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1954_t(x : std_logic_vector) return int1954_t is
  variable rv : int1954_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1955_t_to_slv(x : uint1955_t) return std_logic_vector is
  variable rv : std_logic_vector(1954 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1955_t(x : std_logic_vector) return uint1955_t is
  variable rv : uint1955_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1955_t_to_slv(x : int1955_t) return std_logic_vector is
  variable rv : std_logic_vector(1954 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1955_t(x : std_logic_vector) return int1955_t is
  variable rv : int1955_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1956_t_to_slv(x : uint1956_t) return std_logic_vector is
  variable rv : std_logic_vector(1955 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1956_t(x : std_logic_vector) return uint1956_t is
  variable rv : uint1956_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1956_t_to_slv(x : int1956_t) return std_logic_vector is
  variable rv : std_logic_vector(1955 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1956_t(x : std_logic_vector) return int1956_t is
  variable rv : int1956_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1957_t_to_slv(x : uint1957_t) return std_logic_vector is
  variable rv : std_logic_vector(1956 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1957_t(x : std_logic_vector) return uint1957_t is
  variable rv : uint1957_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1957_t_to_slv(x : int1957_t) return std_logic_vector is
  variable rv : std_logic_vector(1956 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1957_t(x : std_logic_vector) return int1957_t is
  variable rv : int1957_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1958_t_to_slv(x : uint1958_t) return std_logic_vector is
  variable rv : std_logic_vector(1957 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1958_t(x : std_logic_vector) return uint1958_t is
  variable rv : uint1958_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1958_t_to_slv(x : int1958_t) return std_logic_vector is
  variable rv : std_logic_vector(1957 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1958_t(x : std_logic_vector) return int1958_t is
  variable rv : int1958_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1959_t_to_slv(x : uint1959_t) return std_logic_vector is
  variable rv : std_logic_vector(1958 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1959_t(x : std_logic_vector) return uint1959_t is
  variable rv : uint1959_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1959_t_to_slv(x : int1959_t) return std_logic_vector is
  variable rv : std_logic_vector(1958 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1959_t(x : std_logic_vector) return int1959_t is
  variable rv : int1959_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1960_t_to_slv(x : uint1960_t) return std_logic_vector is
  variable rv : std_logic_vector(1959 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1960_t(x : std_logic_vector) return uint1960_t is
  variable rv : uint1960_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1960_t_to_slv(x : int1960_t) return std_logic_vector is
  variable rv : std_logic_vector(1959 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1960_t(x : std_logic_vector) return int1960_t is
  variable rv : int1960_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1961_t_to_slv(x : uint1961_t) return std_logic_vector is
  variable rv : std_logic_vector(1960 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1961_t(x : std_logic_vector) return uint1961_t is
  variable rv : uint1961_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1961_t_to_slv(x : int1961_t) return std_logic_vector is
  variable rv : std_logic_vector(1960 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1961_t(x : std_logic_vector) return int1961_t is
  variable rv : int1961_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1962_t_to_slv(x : uint1962_t) return std_logic_vector is
  variable rv : std_logic_vector(1961 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1962_t(x : std_logic_vector) return uint1962_t is
  variable rv : uint1962_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1962_t_to_slv(x : int1962_t) return std_logic_vector is
  variable rv : std_logic_vector(1961 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1962_t(x : std_logic_vector) return int1962_t is
  variable rv : int1962_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1963_t_to_slv(x : uint1963_t) return std_logic_vector is
  variable rv : std_logic_vector(1962 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1963_t(x : std_logic_vector) return uint1963_t is
  variable rv : uint1963_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1963_t_to_slv(x : int1963_t) return std_logic_vector is
  variable rv : std_logic_vector(1962 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1963_t(x : std_logic_vector) return int1963_t is
  variable rv : int1963_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1964_t_to_slv(x : uint1964_t) return std_logic_vector is
  variable rv : std_logic_vector(1963 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1964_t(x : std_logic_vector) return uint1964_t is
  variable rv : uint1964_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1964_t_to_slv(x : int1964_t) return std_logic_vector is
  variable rv : std_logic_vector(1963 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1964_t(x : std_logic_vector) return int1964_t is
  variable rv : int1964_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1965_t_to_slv(x : uint1965_t) return std_logic_vector is
  variable rv : std_logic_vector(1964 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1965_t(x : std_logic_vector) return uint1965_t is
  variable rv : uint1965_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1965_t_to_slv(x : int1965_t) return std_logic_vector is
  variable rv : std_logic_vector(1964 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1965_t(x : std_logic_vector) return int1965_t is
  variable rv : int1965_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1966_t_to_slv(x : uint1966_t) return std_logic_vector is
  variable rv : std_logic_vector(1965 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1966_t(x : std_logic_vector) return uint1966_t is
  variable rv : uint1966_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1966_t_to_slv(x : int1966_t) return std_logic_vector is
  variable rv : std_logic_vector(1965 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1966_t(x : std_logic_vector) return int1966_t is
  variable rv : int1966_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1967_t_to_slv(x : uint1967_t) return std_logic_vector is
  variable rv : std_logic_vector(1966 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1967_t(x : std_logic_vector) return uint1967_t is
  variable rv : uint1967_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1967_t_to_slv(x : int1967_t) return std_logic_vector is
  variable rv : std_logic_vector(1966 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1967_t(x : std_logic_vector) return int1967_t is
  variable rv : int1967_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1968_t_to_slv(x : uint1968_t) return std_logic_vector is
  variable rv : std_logic_vector(1967 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1968_t(x : std_logic_vector) return uint1968_t is
  variable rv : uint1968_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1968_t_to_slv(x : int1968_t) return std_logic_vector is
  variable rv : std_logic_vector(1967 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1968_t(x : std_logic_vector) return int1968_t is
  variable rv : int1968_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1969_t_to_slv(x : uint1969_t) return std_logic_vector is
  variable rv : std_logic_vector(1968 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1969_t(x : std_logic_vector) return uint1969_t is
  variable rv : uint1969_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1969_t_to_slv(x : int1969_t) return std_logic_vector is
  variable rv : std_logic_vector(1968 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1969_t(x : std_logic_vector) return int1969_t is
  variable rv : int1969_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1970_t_to_slv(x : uint1970_t) return std_logic_vector is
  variable rv : std_logic_vector(1969 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1970_t(x : std_logic_vector) return uint1970_t is
  variable rv : uint1970_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1970_t_to_slv(x : int1970_t) return std_logic_vector is
  variable rv : std_logic_vector(1969 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1970_t(x : std_logic_vector) return int1970_t is
  variable rv : int1970_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1971_t_to_slv(x : uint1971_t) return std_logic_vector is
  variable rv : std_logic_vector(1970 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1971_t(x : std_logic_vector) return uint1971_t is
  variable rv : uint1971_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1971_t_to_slv(x : int1971_t) return std_logic_vector is
  variable rv : std_logic_vector(1970 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1971_t(x : std_logic_vector) return int1971_t is
  variable rv : int1971_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1972_t_to_slv(x : uint1972_t) return std_logic_vector is
  variable rv : std_logic_vector(1971 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1972_t(x : std_logic_vector) return uint1972_t is
  variable rv : uint1972_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1972_t_to_slv(x : int1972_t) return std_logic_vector is
  variable rv : std_logic_vector(1971 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1972_t(x : std_logic_vector) return int1972_t is
  variable rv : int1972_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1973_t_to_slv(x : uint1973_t) return std_logic_vector is
  variable rv : std_logic_vector(1972 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1973_t(x : std_logic_vector) return uint1973_t is
  variable rv : uint1973_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1973_t_to_slv(x : int1973_t) return std_logic_vector is
  variable rv : std_logic_vector(1972 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1973_t(x : std_logic_vector) return int1973_t is
  variable rv : int1973_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1974_t_to_slv(x : uint1974_t) return std_logic_vector is
  variable rv : std_logic_vector(1973 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1974_t(x : std_logic_vector) return uint1974_t is
  variable rv : uint1974_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1974_t_to_slv(x : int1974_t) return std_logic_vector is
  variable rv : std_logic_vector(1973 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1974_t(x : std_logic_vector) return int1974_t is
  variable rv : int1974_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1975_t_to_slv(x : uint1975_t) return std_logic_vector is
  variable rv : std_logic_vector(1974 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1975_t(x : std_logic_vector) return uint1975_t is
  variable rv : uint1975_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1975_t_to_slv(x : int1975_t) return std_logic_vector is
  variable rv : std_logic_vector(1974 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1975_t(x : std_logic_vector) return int1975_t is
  variable rv : int1975_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1976_t_to_slv(x : uint1976_t) return std_logic_vector is
  variable rv : std_logic_vector(1975 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1976_t(x : std_logic_vector) return uint1976_t is
  variable rv : uint1976_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1976_t_to_slv(x : int1976_t) return std_logic_vector is
  variable rv : std_logic_vector(1975 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1976_t(x : std_logic_vector) return int1976_t is
  variable rv : int1976_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1977_t_to_slv(x : uint1977_t) return std_logic_vector is
  variable rv : std_logic_vector(1976 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1977_t(x : std_logic_vector) return uint1977_t is
  variable rv : uint1977_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1977_t_to_slv(x : int1977_t) return std_logic_vector is
  variable rv : std_logic_vector(1976 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1977_t(x : std_logic_vector) return int1977_t is
  variable rv : int1977_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1978_t_to_slv(x : uint1978_t) return std_logic_vector is
  variable rv : std_logic_vector(1977 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1978_t(x : std_logic_vector) return uint1978_t is
  variable rv : uint1978_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1978_t_to_slv(x : int1978_t) return std_logic_vector is
  variable rv : std_logic_vector(1977 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1978_t(x : std_logic_vector) return int1978_t is
  variable rv : int1978_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1979_t_to_slv(x : uint1979_t) return std_logic_vector is
  variable rv : std_logic_vector(1978 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1979_t(x : std_logic_vector) return uint1979_t is
  variable rv : uint1979_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1979_t_to_slv(x : int1979_t) return std_logic_vector is
  variable rv : std_logic_vector(1978 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1979_t(x : std_logic_vector) return int1979_t is
  variable rv : int1979_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1980_t_to_slv(x : uint1980_t) return std_logic_vector is
  variable rv : std_logic_vector(1979 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1980_t(x : std_logic_vector) return uint1980_t is
  variable rv : uint1980_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1980_t_to_slv(x : int1980_t) return std_logic_vector is
  variable rv : std_logic_vector(1979 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1980_t(x : std_logic_vector) return int1980_t is
  variable rv : int1980_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1981_t_to_slv(x : uint1981_t) return std_logic_vector is
  variable rv : std_logic_vector(1980 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1981_t(x : std_logic_vector) return uint1981_t is
  variable rv : uint1981_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1981_t_to_slv(x : int1981_t) return std_logic_vector is
  variable rv : std_logic_vector(1980 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1981_t(x : std_logic_vector) return int1981_t is
  variable rv : int1981_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1982_t_to_slv(x : uint1982_t) return std_logic_vector is
  variable rv : std_logic_vector(1981 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1982_t(x : std_logic_vector) return uint1982_t is
  variable rv : uint1982_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1982_t_to_slv(x : int1982_t) return std_logic_vector is
  variable rv : std_logic_vector(1981 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1982_t(x : std_logic_vector) return int1982_t is
  variable rv : int1982_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1983_t_to_slv(x : uint1983_t) return std_logic_vector is
  variable rv : std_logic_vector(1982 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1983_t(x : std_logic_vector) return uint1983_t is
  variable rv : uint1983_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1983_t_to_slv(x : int1983_t) return std_logic_vector is
  variable rv : std_logic_vector(1982 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1983_t(x : std_logic_vector) return int1983_t is
  variable rv : int1983_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1984_t_to_slv(x : uint1984_t) return std_logic_vector is
  variable rv : std_logic_vector(1983 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1984_t(x : std_logic_vector) return uint1984_t is
  variable rv : uint1984_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1984_t_to_slv(x : int1984_t) return std_logic_vector is
  variable rv : std_logic_vector(1983 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1984_t(x : std_logic_vector) return int1984_t is
  variable rv : int1984_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1985_t_to_slv(x : uint1985_t) return std_logic_vector is
  variable rv : std_logic_vector(1984 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1985_t(x : std_logic_vector) return uint1985_t is
  variable rv : uint1985_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1985_t_to_slv(x : int1985_t) return std_logic_vector is
  variable rv : std_logic_vector(1984 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1985_t(x : std_logic_vector) return int1985_t is
  variable rv : int1985_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1986_t_to_slv(x : uint1986_t) return std_logic_vector is
  variable rv : std_logic_vector(1985 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1986_t(x : std_logic_vector) return uint1986_t is
  variable rv : uint1986_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1986_t_to_slv(x : int1986_t) return std_logic_vector is
  variable rv : std_logic_vector(1985 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1986_t(x : std_logic_vector) return int1986_t is
  variable rv : int1986_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1987_t_to_slv(x : uint1987_t) return std_logic_vector is
  variable rv : std_logic_vector(1986 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1987_t(x : std_logic_vector) return uint1987_t is
  variable rv : uint1987_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1987_t_to_slv(x : int1987_t) return std_logic_vector is
  variable rv : std_logic_vector(1986 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1987_t(x : std_logic_vector) return int1987_t is
  variable rv : int1987_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1988_t_to_slv(x : uint1988_t) return std_logic_vector is
  variable rv : std_logic_vector(1987 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1988_t(x : std_logic_vector) return uint1988_t is
  variable rv : uint1988_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1988_t_to_slv(x : int1988_t) return std_logic_vector is
  variable rv : std_logic_vector(1987 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1988_t(x : std_logic_vector) return int1988_t is
  variable rv : int1988_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1989_t_to_slv(x : uint1989_t) return std_logic_vector is
  variable rv : std_logic_vector(1988 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1989_t(x : std_logic_vector) return uint1989_t is
  variable rv : uint1989_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1989_t_to_slv(x : int1989_t) return std_logic_vector is
  variable rv : std_logic_vector(1988 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1989_t(x : std_logic_vector) return int1989_t is
  variable rv : int1989_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1990_t_to_slv(x : uint1990_t) return std_logic_vector is
  variable rv : std_logic_vector(1989 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1990_t(x : std_logic_vector) return uint1990_t is
  variable rv : uint1990_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1990_t_to_slv(x : int1990_t) return std_logic_vector is
  variable rv : std_logic_vector(1989 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1990_t(x : std_logic_vector) return int1990_t is
  variable rv : int1990_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1991_t_to_slv(x : uint1991_t) return std_logic_vector is
  variable rv : std_logic_vector(1990 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1991_t(x : std_logic_vector) return uint1991_t is
  variable rv : uint1991_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1991_t_to_slv(x : int1991_t) return std_logic_vector is
  variable rv : std_logic_vector(1990 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1991_t(x : std_logic_vector) return int1991_t is
  variable rv : int1991_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1992_t_to_slv(x : uint1992_t) return std_logic_vector is
  variable rv : std_logic_vector(1991 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1992_t(x : std_logic_vector) return uint1992_t is
  variable rv : uint1992_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1992_t_to_slv(x : int1992_t) return std_logic_vector is
  variable rv : std_logic_vector(1991 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1992_t(x : std_logic_vector) return int1992_t is
  variable rv : int1992_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1993_t_to_slv(x : uint1993_t) return std_logic_vector is
  variable rv : std_logic_vector(1992 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1993_t(x : std_logic_vector) return uint1993_t is
  variable rv : uint1993_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1993_t_to_slv(x : int1993_t) return std_logic_vector is
  variable rv : std_logic_vector(1992 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1993_t(x : std_logic_vector) return int1993_t is
  variable rv : int1993_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1994_t_to_slv(x : uint1994_t) return std_logic_vector is
  variable rv : std_logic_vector(1993 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1994_t(x : std_logic_vector) return uint1994_t is
  variable rv : uint1994_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1994_t_to_slv(x : int1994_t) return std_logic_vector is
  variable rv : std_logic_vector(1993 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1994_t(x : std_logic_vector) return int1994_t is
  variable rv : int1994_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1995_t_to_slv(x : uint1995_t) return std_logic_vector is
  variable rv : std_logic_vector(1994 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1995_t(x : std_logic_vector) return uint1995_t is
  variable rv : uint1995_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1995_t_to_slv(x : int1995_t) return std_logic_vector is
  variable rv : std_logic_vector(1994 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1995_t(x : std_logic_vector) return int1995_t is
  variable rv : int1995_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1996_t_to_slv(x : uint1996_t) return std_logic_vector is
  variable rv : std_logic_vector(1995 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1996_t(x : std_logic_vector) return uint1996_t is
  variable rv : uint1996_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1996_t_to_slv(x : int1996_t) return std_logic_vector is
  variable rv : std_logic_vector(1995 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1996_t(x : std_logic_vector) return int1996_t is
  variable rv : int1996_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1997_t_to_slv(x : uint1997_t) return std_logic_vector is
  variable rv : std_logic_vector(1996 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1997_t(x : std_logic_vector) return uint1997_t is
  variable rv : uint1997_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1997_t_to_slv(x : int1997_t) return std_logic_vector is
  variable rv : std_logic_vector(1996 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1997_t(x : std_logic_vector) return int1997_t is
  variable rv : int1997_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1998_t_to_slv(x : uint1998_t) return std_logic_vector is
  variable rv : std_logic_vector(1997 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1998_t(x : std_logic_vector) return uint1998_t is
  variable rv : uint1998_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1998_t_to_slv(x : int1998_t) return std_logic_vector is
  variable rv : std_logic_vector(1997 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1998_t(x : std_logic_vector) return int1998_t is
  variable rv : int1998_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint1999_t_to_slv(x : uint1999_t) return std_logic_vector is
  variable rv : std_logic_vector(1998 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint1999_t(x : std_logic_vector) return uint1999_t is
  variable rv : uint1999_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int1999_t_to_slv(x : int1999_t) return std_logic_vector is
  variable rv : std_logic_vector(1998 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int1999_t(x : std_logic_vector) return int1999_t is
  variable rv : int1999_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2000_t_to_slv(x : uint2000_t) return std_logic_vector is
  variable rv : std_logic_vector(1999 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2000_t(x : std_logic_vector) return uint2000_t is
  variable rv : uint2000_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2000_t_to_slv(x : int2000_t) return std_logic_vector is
  variable rv : std_logic_vector(1999 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2000_t(x : std_logic_vector) return int2000_t is
  variable rv : int2000_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2001_t_to_slv(x : uint2001_t) return std_logic_vector is
  variable rv : std_logic_vector(2000 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2001_t(x : std_logic_vector) return uint2001_t is
  variable rv : uint2001_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2001_t_to_slv(x : int2001_t) return std_logic_vector is
  variable rv : std_logic_vector(2000 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2001_t(x : std_logic_vector) return int2001_t is
  variable rv : int2001_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2002_t_to_slv(x : uint2002_t) return std_logic_vector is
  variable rv : std_logic_vector(2001 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2002_t(x : std_logic_vector) return uint2002_t is
  variable rv : uint2002_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2002_t_to_slv(x : int2002_t) return std_logic_vector is
  variable rv : std_logic_vector(2001 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2002_t(x : std_logic_vector) return int2002_t is
  variable rv : int2002_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2003_t_to_slv(x : uint2003_t) return std_logic_vector is
  variable rv : std_logic_vector(2002 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2003_t(x : std_logic_vector) return uint2003_t is
  variable rv : uint2003_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2003_t_to_slv(x : int2003_t) return std_logic_vector is
  variable rv : std_logic_vector(2002 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2003_t(x : std_logic_vector) return int2003_t is
  variable rv : int2003_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2004_t_to_slv(x : uint2004_t) return std_logic_vector is
  variable rv : std_logic_vector(2003 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2004_t(x : std_logic_vector) return uint2004_t is
  variable rv : uint2004_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2004_t_to_slv(x : int2004_t) return std_logic_vector is
  variable rv : std_logic_vector(2003 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2004_t(x : std_logic_vector) return int2004_t is
  variable rv : int2004_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2005_t_to_slv(x : uint2005_t) return std_logic_vector is
  variable rv : std_logic_vector(2004 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2005_t(x : std_logic_vector) return uint2005_t is
  variable rv : uint2005_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2005_t_to_slv(x : int2005_t) return std_logic_vector is
  variable rv : std_logic_vector(2004 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2005_t(x : std_logic_vector) return int2005_t is
  variable rv : int2005_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2006_t_to_slv(x : uint2006_t) return std_logic_vector is
  variable rv : std_logic_vector(2005 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2006_t(x : std_logic_vector) return uint2006_t is
  variable rv : uint2006_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2006_t_to_slv(x : int2006_t) return std_logic_vector is
  variable rv : std_logic_vector(2005 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2006_t(x : std_logic_vector) return int2006_t is
  variable rv : int2006_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2007_t_to_slv(x : uint2007_t) return std_logic_vector is
  variable rv : std_logic_vector(2006 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2007_t(x : std_logic_vector) return uint2007_t is
  variable rv : uint2007_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2007_t_to_slv(x : int2007_t) return std_logic_vector is
  variable rv : std_logic_vector(2006 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2007_t(x : std_logic_vector) return int2007_t is
  variable rv : int2007_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2008_t_to_slv(x : uint2008_t) return std_logic_vector is
  variable rv : std_logic_vector(2007 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2008_t(x : std_logic_vector) return uint2008_t is
  variable rv : uint2008_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2008_t_to_slv(x : int2008_t) return std_logic_vector is
  variable rv : std_logic_vector(2007 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2008_t(x : std_logic_vector) return int2008_t is
  variable rv : int2008_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2009_t_to_slv(x : uint2009_t) return std_logic_vector is
  variable rv : std_logic_vector(2008 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2009_t(x : std_logic_vector) return uint2009_t is
  variable rv : uint2009_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2009_t_to_slv(x : int2009_t) return std_logic_vector is
  variable rv : std_logic_vector(2008 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2009_t(x : std_logic_vector) return int2009_t is
  variable rv : int2009_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2010_t_to_slv(x : uint2010_t) return std_logic_vector is
  variable rv : std_logic_vector(2009 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2010_t(x : std_logic_vector) return uint2010_t is
  variable rv : uint2010_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2010_t_to_slv(x : int2010_t) return std_logic_vector is
  variable rv : std_logic_vector(2009 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2010_t(x : std_logic_vector) return int2010_t is
  variable rv : int2010_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2011_t_to_slv(x : uint2011_t) return std_logic_vector is
  variable rv : std_logic_vector(2010 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2011_t(x : std_logic_vector) return uint2011_t is
  variable rv : uint2011_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2011_t_to_slv(x : int2011_t) return std_logic_vector is
  variable rv : std_logic_vector(2010 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2011_t(x : std_logic_vector) return int2011_t is
  variable rv : int2011_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2012_t_to_slv(x : uint2012_t) return std_logic_vector is
  variable rv : std_logic_vector(2011 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2012_t(x : std_logic_vector) return uint2012_t is
  variable rv : uint2012_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2012_t_to_slv(x : int2012_t) return std_logic_vector is
  variable rv : std_logic_vector(2011 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2012_t(x : std_logic_vector) return int2012_t is
  variable rv : int2012_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2013_t_to_slv(x : uint2013_t) return std_logic_vector is
  variable rv : std_logic_vector(2012 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2013_t(x : std_logic_vector) return uint2013_t is
  variable rv : uint2013_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2013_t_to_slv(x : int2013_t) return std_logic_vector is
  variable rv : std_logic_vector(2012 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2013_t(x : std_logic_vector) return int2013_t is
  variable rv : int2013_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2014_t_to_slv(x : uint2014_t) return std_logic_vector is
  variable rv : std_logic_vector(2013 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2014_t(x : std_logic_vector) return uint2014_t is
  variable rv : uint2014_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2014_t_to_slv(x : int2014_t) return std_logic_vector is
  variable rv : std_logic_vector(2013 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2014_t(x : std_logic_vector) return int2014_t is
  variable rv : int2014_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2015_t_to_slv(x : uint2015_t) return std_logic_vector is
  variable rv : std_logic_vector(2014 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2015_t(x : std_logic_vector) return uint2015_t is
  variable rv : uint2015_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2015_t_to_slv(x : int2015_t) return std_logic_vector is
  variable rv : std_logic_vector(2014 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2015_t(x : std_logic_vector) return int2015_t is
  variable rv : int2015_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2016_t_to_slv(x : uint2016_t) return std_logic_vector is
  variable rv : std_logic_vector(2015 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2016_t(x : std_logic_vector) return uint2016_t is
  variable rv : uint2016_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2016_t_to_slv(x : int2016_t) return std_logic_vector is
  variable rv : std_logic_vector(2015 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2016_t(x : std_logic_vector) return int2016_t is
  variable rv : int2016_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2017_t_to_slv(x : uint2017_t) return std_logic_vector is
  variable rv : std_logic_vector(2016 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2017_t(x : std_logic_vector) return uint2017_t is
  variable rv : uint2017_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2017_t_to_slv(x : int2017_t) return std_logic_vector is
  variable rv : std_logic_vector(2016 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2017_t(x : std_logic_vector) return int2017_t is
  variable rv : int2017_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2018_t_to_slv(x : uint2018_t) return std_logic_vector is
  variable rv : std_logic_vector(2017 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2018_t(x : std_logic_vector) return uint2018_t is
  variable rv : uint2018_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2018_t_to_slv(x : int2018_t) return std_logic_vector is
  variable rv : std_logic_vector(2017 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2018_t(x : std_logic_vector) return int2018_t is
  variable rv : int2018_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2019_t_to_slv(x : uint2019_t) return std_logic_vector is
  variable rv : std_logic_vector(2018 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2019_t(x : std_logic_vector) return uint2019_t is
  variable rv : uint2019_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2019_t_to_slv(x : int2019_t) return std_logic_vector is
  variable rv : std_logic_vector(2018 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2019_t(x : std_logic_vector) return int2019_t is
  variable rv : int2019_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2020_t_to_slv(x : uint2020_t) return std_logic_vector is
  variable rv : std_logic_vector(2019 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2020_t(x : std_logic_vector) return uint2020_t is
  variable rv : uint2020_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2020_t_to_slv(x : int2020_t) return std_logic_vector is
  variable rv : std_logic_vector(2019 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2020_t(x : std_logic_vector) return int2020_t is
  variable rv : int2020_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2021_t_to_slv(x : uint2021_t) return std_logic_vector is
  variable rv : std_logic_vector(2020 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2021_t(x : std_logic_vector) return uint2021_t is
  variable rv : uint2021_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2021_t_to_slv(x : int2021_t) return std_logic_vector is
  variable rv : std_logic_vector(2020 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2021_t(x : std_logic_vector) return int2021_t is
  variable rv : int2021_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2022_t_to_slv(x : uint2022_t) return std_logic_vector is
  variable rv : std_logic_vector(2021 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2022_t(x : std_logic_vector) return uint2022_t is
  variable rv : uint2022_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2022_t_to_slv(x : int2022_t) return std_logic_vector is
  variable rv : std_logic_vector(2021 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2022_t(x : std_logic_vector) return int2022_t is
  variable rv : int2022_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2023_t_to_slv(x : uint2023_t) return std_logic_vector is
  variable rv : std_logic_vector(2022 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2023_t(x : std_logic_vector) return uint2023_t is
  variable rv : uint2023_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2023_t_to_slv(x : int2023_t) return std_logic_vector is
  variable rv : std_logic_vector(2022 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2023_t(x : std_logic_vector) return int2023_t is
  variable rv : int2023_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2024_t_to_slv(x : uint2024_t) return std_logic_vector is
  variable rv : std_logic_vector(2023 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2024_t(x : std_logic_vector) return uint2024_t is
  variable rv : uint2024_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2024_t_to_slv(x : int2024_t) return std_logic_vector is
  variable rv : std_logic_vector(2023 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2024_t(x : std_logic_vector) return int2024_t is
  variable rv : int2024_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2025_t_to_slv(x : uint2025_t) return std_logic_vector is
  variable rv : std_logic_vector(2024 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2025_t(x : std_logic_vector) return uint2025_t is
  variable rv : uint2025_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2025_t_to_slv(x : int2025_t) return std_logic_vector is
  variable rv : std_logic_vector(2024 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2025_t(x : std_logic_vector) return int2025_t is
  variable rv : int2025_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2026_t_to_slv(x : uint2026_t) return std_logic_vector is
  variable rv : std_logic_vector(2025 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2026_t(x : std_logic_vector) return uint2026_t is
  variable rv : uint2026_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2026_t_to_slv(x : int2026_t) return std_logic_vector is
  variable rv : std_logic_vector(2025 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2026_t(x : std_logic_vector) return int2026_t is
  variable rv : int2026_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2027_t_to_slv(x : uint2027_t) return std_logic_vector is
  variable rv : std_logic_vector(2026 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2027_t(x : std_logic_vector) return uint2027_t is
  variable rv : uint2027_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2027_t_to_slv(x : int2027_t) return std_logic_vector is
  variable rv : std_logic_vector(2026 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2027_t(x : std_logic_vector) return int2027_t is
  variable rv : int2027_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2028_t_to_slv(x : uint2028_t) return std_logic_vector is
  variable rv : std_logic_vector(2027 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2028_t(x : std_logic_vector) return uint2028_t is
  variable rv : uint2028_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2028_t_to_slv(x : int2028_t) return std_logic_vector is
  variable rv : std_logic_vector(2027 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2028_t(x : std_logic_vector) return int2028_t is
  variable rv : int2028_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2029_t_to_slv(x : uint2029_t) return std_logic_vector is
  variable rv : std_logic_vector(2028 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2029_t(x : std_logic_vector) return uint2029_t is
  variable rv : uint2029_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2029_t_to_slv(x : int2029_t) return std_logic_vector is
  variable rv : std_logic_vector(2028 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2029_t(x : std_logic_vector) return int2029_t is
  variable rv : int2029_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2030_t_to_slv(x : uint2030_t) return std_logic_vector is
  variable rv : std_logic_vector(2029 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2030_t(x : std_logic_vector) return uint2030_t is
  variable rv : uint2030_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2030_t_to_slv(x : int2030_t) return std_logic_vector is
  variable rv : std_logic_vector(2029 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2030_t(x : std_logic_vector) return int2030_t is
  variable rv : int2030_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2031_t_to_slv(x : uint2031_t) return std_logic_vector is
  variable rv : std_logic_vector(2030 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2031_t(x : std_logic_vector) return uint2031_t is
  variable rv : uint2031_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2031_t_to_slv(x : int2031_t) return std_logic_vector is
  variable rv : std_logic_vector(2030 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2031_t(x : std_logic_vector) return int2031_t is
  variable rv : int2031_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2032_t_to_slv(x : uint2032_t) return std_logic_vector is
  variable rv : std_logic_vector(2031 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2032_t(x : std_logic_vector) return uint2032_t is
  variable rv : uint2032_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2032_t_to_slv(x : int2032_t) return std_logic_vector is
  variable rv : std_logic_vector(2031 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2032_t(x : std_logic_vector) return int2032_t is
  variable rv : int2032_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2033_t_to_slv(x : uint2033_t) return std_logic_vector is
  variable rv : std_logic_vector(2032 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2033_t(x : std_logic_vector) return uint2033_t is
  variable rv : uint2033_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2033_t_to_slv(x : int2033_t) return std_logic_vector is
  variable rv : std_logic_vector(2032 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2033_t(x : std_logic_vector) return int2033_t is
  variable rv : int2033_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2034_t_to_slv(x : uint2034_t) return std_logic_vector is
  variable rv : std_logic_vector(2033 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2034_t(x : std_logic_vector) return uint2034_t is
  variable rv : uint2034_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2034_t_to_slv(x : int2034_t) return std_logic_vector is
  variable rv : std_logic_vector(2033 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2034_t(x : std_logic_vector) return int2034_t is
  variable rv : int2034_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2035_t_to_slv(x : uint2035_t) return std_logic_vector is
  variable rv : std_logic_vector(2034 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2035_t(x : std_logic_vector) return uint2035_t is
  variable rv : uint2035_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2035_t_to_slv(x : int2035_t) return std_logic_vector is
  variable rv : std_logic_vector(2034 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2035_t(x : std_logic_vector) return int2035_t is
  variable rv : int2035_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2036_t_to_slv(x : uint2036_t) return std_logic_vector is
  variable rv : std_logic_vector(2035 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2036_t(x : std_logic_vector) return uint2036_t is
  variable rv : uint2036_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2036_t_to_slv(x : int2036_t) return std_logic_vector is
  variable rv : std_logic_vector(2035 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2036_t(x : std_logic_vector) return int2036_t is
  variable rv : int2036_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2037_t_to_slv(x : uint2037_t) return std_logic_vector is
  variable rv : std_logic_vector(2036 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2037_t(x : std_logic_vector) return uint2037_t is
  variable rv : uint2037_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2037_t_to_slv(x : int2037_t) return std_logic_vector is
  variable rv : std_logic_vector(2036 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2037_t(x : std_logic_vector) return int2037_t is
  variable rv : int2037_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2038_t_to_slv(x : uint2038_t) return std_logic_vector is
  variable rv : std_logic_vector(2037 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2038_t(x : std_logic_vector) return uint2038_t is
  variable rv : uint2038_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2038_t_to_slv(x : int2038_t) return std_logic_vector is
  variable rv : std_logic_vector(2037 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2038_t(x : std_logic_vector) return int2038_t is
  variable rv : int2038_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2039_t_to_slv(x : uint2039_t) return std_logic_vector is
  variable rv : std_logic_vector(2038 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2039_t(x : std_logic_vector) return uint2039_t is
  variable rv : uint2039_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2039_t_to_slv(x : int2039_t) return std_logic_vector is
  variable rv : std_logic_vector(2038 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2039_t(x : std_logic_vector) return int2039_t is
  variable rv : int2039_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2040_t_to_slv(x : uint2040_t) return std_logic_vector is
  variable rv : std_logic_vector(2039 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2040_t(x : std_logic_vector) return uint2040_t is
  variable rv : uint2040_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2040_t_to_slv(x : int2040_t) return std_logic_vector is
  variable rv : std_logic_vector(2039 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2040_t(x : std_logic_vector) return int2040_t is
  variable rv : int2040_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2041_t_to_slv(x : uint2041_t) return std_logic_vector is
  variable rv : std_logic_vector(2040 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2041_t(x : std_logic_vector) return uint2041_t is
  variable rv : uint2041_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2041_t_to_slv(x : int2041_t) return std_logic_vector is
  variable rv : std_logic_vector(2040 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2041_t(x : std_logic_vector) return int2041_t is
  variable rv : int2041_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2042_t_to_slv(x : uint2042_t) return std_logic_vector is
  variable rv : std_logic_vector(2041 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2042_t(x : std_logic_vector) return uint2042_t is
  variable rv : uint2042_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2042_t_to_slv(x : int2042_t) return std_logic_vector is
  variable rv : std_logic_vector(2041 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2042_t(x : std_logic_vector) return int2042_t is
  variable rv : int2042_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2043_t_to_slv(x : uint2043_t) return std_logic_vector is
  variable rv : std_logic_vector(2042 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2043_t(x : std_logic_vector) return uint2043_t is
  variable rv : uint2043_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2043_t_to_slv(x : int2043_t) return std_logic_vector is
  variable rv : std_logic_vector(2042 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2043_t(x : std_logic_vector) return int2043_t is
  variable rv : int2043_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2044_t_to_slv(x : uint2044_t) return std_logic_vector is
  variable rv : std_logic_vector(2043 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2044_t(x : std_logic_vector) return uint2044_t is
  variable rv : uint2044_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2044_t_to_slv(x : int2044_t) return std_logic_vector is
  variable rv : std_logic_vector(2043 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2044_t(x : std_logic_vector) return int2044_t is
  variable rv : int2044_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2045_t_to_slv(x : uint2045_t) return std_logic_vector is
  variable rv : std_logic_vector(2044 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2045_t(x : std_logic_vector) return uint2045_t is
  variable rv : uint2045_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2045_t_to_slv(x : int2045_t) return std_logic_vector is
  variable rv : std_logic_vector(2044 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2045_t(x : std_logic_vector) return int2045_t is
  variable rv : int2045_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2046_t_to_slv(x : uint2046_t) return std_logic_vector is
  variable rv : std_logic_vector(2045 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2046_t(x : std_logic_vector) return uint2046_t is
  variable rv : uint2046_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2046_t_to_slv(x : int2046_t) return std_logic_vector is
  variable rv : std_logic_vector(2045 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2046_t(x : std_logic_vector) return int2046_t is
  variable rv : int2046_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2047_t_to_slv(x : uint2047_t) return std_logic_vector is
  variable rv : std_logic_vector(2046 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2047_t(x : std_logic_vector) return uint2047_t is
  variable rv : uint2047_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2047_t_to_slv(x : int2047_t) return std_logic_vector is
  variable rv : std_logic_vector(2046 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2047_t(x : std_logic_vector) return int2047_t is
  variable rv : int2047_t;
begin
    rv := signed(x);
    return rv;
end function;
function uint2048_t_to_slv(x : uint2048_t) return std_logic_vector is
  variable rv : std_logic_vector(2047 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_uint2048_t(x : std_logic_vector) return uint2048_t is
  variable rv : uint2048_t;
begin
    rv := unsigned(x);
    return rv;
end function;
function int2048_t_to_slv(x : int2048_t) return std_logic_vector is
  variable rv : std_logic_vector(2047 downto 0);
begin
  rv := std_logic_vector(x);
  return rv;
end function;
function slv_to_int2048_t(x : std_logic_vector) return int2048_t is
  variable rv : int2048_t;
begin
    rv := signed(x);
    return rv;
end function;

  function to_byte_array(s : string; constant len : natural) return byte_array_t is
    variable rv : byte_array_t(0 to len-1) := (others=> (others=>'0'));
  begin
    for i in 0 to s'length-1 loop
        -- i+1 since strings start at index 1
        rv(i) := to_unsigned(character'pos(s(i+1)), 8);
    end loop;
    return rv;
  end function;
  
  function resize_float_e_m_t(
    x : std_logic_vector; 
    in_exponent_width : integer;
    in_mantissa_width : integer;
    out_exponent_width : integer;
    out_mantissa_width : integer) return std_logic_vector
  is
    variable x_s : std_logic;
    variable x_e : signed(in_exponent_width-1 downto 0);
    variable x_m : unsigned(in_mantissa_width-1 downto 0);
    variable x_bias : integer := (2**(in_exponent_width-1)) - 1;
    variable rv_s : std_logic;
    variable rv_e : signed(out_exponent_width-1 downto 0);
    variable rv_m : unsigned(out_mantissa_width-1 downto 0);
    variable rv_bias : integer := (2**(out_exponent_width-1)) - 1;
    variable rv : std_logic_vector((1+out_exponent_width+out_mantissa_width)-1 downto 0);
  begin
    x_s := x(in_exponent_width+in_mantissa_width);
    x_e := signed(x((in_exponent_width+in_mantissa_width)-1 downto in_mantissa_width));
    x_m := unsigned(x(in_mantissa_width-1 downto 0));
    
    -- Default zero
    rv_s := x_s;
    rv_e := (others => '0');
    rv_m := (others => '0');
    
    -- Check if non zero
    if not(x_e = to_signed(0, in_exponent_width)) then
      -- Exponent change bias
      rv_e := resize(signed('0' & x_e) - x_bias, out_exponent_width); -- De-bias
      rv_e := rv_e + rv_bias; -- Re-bias
            
      -- Top left n bits of mantissa
      if out_mantissa_width <= in_mantissa_width then
        rv_m := x_m(in_mantissa_width-1 downto (in_mantissa_width-out_mantissa_width));
      else
        -- All bits padded with zeros on right
        rv_m := x_m & to_unsigned(0, out_mantissa_width-in_mantissa_width);
      end if;
    end if;
    
    rv := rv_s & std_logic_vector(rv_e) & std_logic_vector(rv_m);
    return rv;
  end function;
function chacha20_decrypt_state_t_to_slv(e : chacha20_decrypt_state_t) return std_logic_vector is
    variable rv: std_logic_vector(0 downto 0) := (others => '0');
begin
case(e) is
when POLY_KEY => rv := std_logic_vector(to_unsigned(0, 1));
when PLAINTEXT => rv := std_logic_vector(to_unsigned(1, 1));

end case;
return rv;
end function;
    
function prep_auth_data_state_t_to_slv(e : prep_auth_data_state_t) return std_logic_vector is
    variable rv: std_logic_vector(1 downto 0) := (others => '0');
begin
case(e) is
when IDLE => rv := std_logic_vector(to_unsigned(0, 2));
when AAD => rv := std_logic_vector(to_unsigned(1, 2));
when CIPHERTEXT => rv := std_logic_vector(to_unsigned(2, 2));
when LENGTHS => rv := std_logic_vector(to_unsigned(3, 2));

end case;
return rv;
end function;
    
function poly1305_state_t_to_slv(e : poly1305_state_t) return std_logic_vector is
    variable rv: std_logic_vector(2 downto 0) := (others => '0');
begin
case(e) is
when IDLE => rv := std_logic_vector(to_unsigned(0, 3));
when START_ITER => rv := std_logic_vector(to_unsigned(1, 3));
when FINISH_ITER => rv := std_logic_vector(to_unsigned(2, 3));
when A_PLUS_S => rv := std_logic_vector(to_unsigned(3, 3));
when OUTPUT_AUTH_TAG => rv := std_logic_vector(to_unsigned(4, 3));

end case;
return rv;
end function;
    
function poly1305_verify_state_t_to_slv(e : poly1305_verify_state_t) return std_logic_vector is
    variable rv: std_logic_vector(1 downto 0) := (others => '0');
begin
case(e) is
when TAKE_AUTH_TAG => rv := std_logic_vector(to_unsigned(0, 2));
when TAKE_CALC_TAG => rv := std_logic_vector(to_unsigned(1, 2));
when COMPARE_TAGS => rv := std_logic_vector(to_unsigned(2, 2));
when OUTPUT_COMPARE_RESULT => rv := std_logic_vector(to_unsigned(3, 2));

end case;
return rv;
end function;
    
function strip_auth_tag_state_t_to_slv(e : strip_auth_tag_state_t) return std_logic_vector is
    variable rv: std_logic_vector(0 downto 0) := (others => '0');
begin
case(e) is
when CIPHERTEXT_PASS => rv := std_logic_vector(to_unsigned(0, 1));
when AUTH_TAG_EXTRACTION => rv := std_logic_vector(to_unsigned(1, 1));

end case;
return rv;
end function;
    
function wait_to_verify_state_t_to_slv(e : wait_to_verify_state_t) return std_logic_vector is
    variable rv: std_logic_vector(0 downto 0) := (others => '0');
begin
case(e) is
when WAIT_TO_VERIFY_BIT => rv := std_logic_vector(to_unsigned(0, 1));
when OUTPUT_PLAINTEXT => rv := std_logic_vector(to_unsigned(1, 1));

end case;
return rv;
end function;
    
      function uint8_t_16_to_slv(data : uint8_t_16) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_16_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_16(data : std_logic_vector) return uint8_t_16 is
        variable rv : uint8_t_16;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function uint64_t_5_to_slv(data : uint64_t_5) return std_logic_vector is
        variable rv : std_logic_vector(uint64_t_5_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+64)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 64;
    
            rv((pos+64)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 64;
    
            rv((pos+64)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 64;
    
            rv((pos+64)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 64;
    
            rv((pos+64)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 64;
    
          return rv;
      end function;
    
      function slv_to_uint64_t_5(data : std_logic_vector) return uint64_t_5 is
        variable rv : uint64_t_5;
        variable elem_slv : std_logic_vector(64-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+64)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 64;
    
            elem_slv := data((pos+64)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 64;
    
            elem_slv := data((pos+64)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 64;
    
            elem_slv := data((pos+64)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 64;
    
            elem_slv := data((pos+64)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 64;
    
          return rv;
      end function;
    
      function uint8_t_32_to_slv(data : uint8_t_32) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_32_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(16));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(17));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(18));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(19));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(20));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(21));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(22));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(23));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(24));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(25));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(26));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(27));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(28));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(29));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(30));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(31));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_32(data : std_logic_vector) return uint8_t_32 is
        variable rv : uint8_t_32;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(16) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(17) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(18) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(19) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(20) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(21) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(22) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(23) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(24) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(25) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(26) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(27) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(28) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(29) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(30) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(31) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function uint8_t_12_to_slv(data : uint8_t_12) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_12_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_12(data : std_logic_vector) return uint8_t_12 is
        variable rv : uint8_t_12;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function uint1_t_64_to_slv(data : uint1_t_64) return std_logic_vector is
        variable rv : std_logic_vector(uint1_t_64_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(16));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(17));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(18));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(19));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(20));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(21));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(22));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(23));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(24));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(25));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(26));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(27));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(28));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(29));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(30));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(31));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(32));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(33));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(34));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(35));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(36));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(37));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(38));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(39));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(40));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(41));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(42));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(43));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(44));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(45));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(46));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(47));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(48));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(49));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(50));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(51));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(52));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(53));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(54));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(55));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(56));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(57));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(58));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(59));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(60));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(61));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(62));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(63));
            pos := pos + 1;
    
          return rv;
      end function;
    
      function slv_to_uint1_t_64(data : std_logic_vector) return uint1_t_64 is
        variable rv : uint1_t_64;
        variable elem_slv : std_logic_vector(1-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(16) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(17) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(18) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(19) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(20) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(21) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(22) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(23) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(24) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(25) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(26) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(27) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(28) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(29) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(30) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(31) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(32) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(33) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(34) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(35) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(36) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(37) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(38) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(39) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(40) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(41) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(42) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(43) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(44) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(45) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(46) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(47) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(48) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(49) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(50) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(51) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(52) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(53) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(54) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(55) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(56) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(57) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(58) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(59) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(60) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(61) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(62) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(63) := unsigned(elem_slv);
            pos := pos + 1;
    
          return rv;
      end function;
    
      function uint1_t_16_to_slv(data : uint1_t_16) return std_logic_vector is
        variable rv : std_logic_vector(uint1_t_16_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 1;
    
          return rv;
      end function;
    
      function slv_to_uint1_t_16(data : std_logic_vector) return uint1_t_16 is
        variable rv : uint1_t_16;
        variable elem_slv : std_logic_vector(1-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 1;
    
          return rv;
      end function;
    
      function uint32_t_8_to_slv(data : uint32_t_8) return std_logic_vector is
        variable rv : std_logic_vector(uint32_t_8_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 32;
    
          return rv;
      end function;
    
      function slv_to_uint32_t_8(data : std_logic_vector) return uint32_t_8 is
        variable rv : uint32_t_8;
        variable elem_slv : std_logic_vector(32-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 32;
    
          return rv;
      end function;
    
      function uint32_t_3_to_slv(data : uint32_t_3) return std_logic_vector is
        variable rv : std_logic_vector(uint32_t_3_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 32;
    
          return rv;
      end function;
    
      function slv_to_uint32_t_3(data : std_logic_vector) return uint32_t_3 is
        variable rv : uint32_t_3;
        variable elem_slv : std_logic_vector(32-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 32;
    
          return rv;
      end function;
    
      function uint8_t_64_to_slv(data : uint8_t_64) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_64_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(16));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(17));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(18));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(19));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(20));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(21));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(22));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(23));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(24));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(25));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(26));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(27));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(28));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(29));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(30));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(31));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(32));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(33));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(34));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(35));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(36));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(37));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(38));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(39));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(40));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(41));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(42));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(43));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(44));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(45));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(46));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(47));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(48));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(49));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(50));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(51));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(52));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(53));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(54));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(55));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(56));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(57));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(58));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(59));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(60));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(61));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(62));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(63));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_64(data : std_logic_vector) return uint8_t_64 is
        variable rv : uint8_t_64;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(16) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(17) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(18) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(19) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(20) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(21) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(22) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(23) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(24) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(25) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(26) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(27) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(28) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(29) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(30) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(31) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(32) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(33) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(34) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(35) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(36) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(37) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(38) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(39) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(40) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(41) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(42) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(43) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(44) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(45) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(46) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(47) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(48) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(49) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(50) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(51) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(52) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(53) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(54) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(55) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(56) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(57) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(58) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(59) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(60) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(61) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(62) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(63) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function uint8_t_8_to_slv(data : uint8_t_8) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_8_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_8(data : std_logic_vector) return uint8_t_8 is
        variable rv : uint8_t_8;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function uint8_t_40_to_slv(data : uint8_t_40) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_40_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(16));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(17));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(18));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(19));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(20));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(21));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(22));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(23));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(24));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(25));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(26));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(27));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(28));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(29));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(30));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(31));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(32));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(33));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(34));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(35));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(36));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(37));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(38));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(39));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_40(data : std_logic_vector) return uint8_t_40 is
        variable rv : uint8_t_40;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(16) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(17) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(18) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(19) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(20) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(21) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(22) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(23) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(24) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(25) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(26) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(27) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(28) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(29) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(30) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(31) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(32) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(33) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(34) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(35) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(36) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(37) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(38) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(39) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function char_128_to_slv(data : char_128) return std_logic_vector is
        variable rv : std_logic_vector(char_128_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(16));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(17));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(18));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(19));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(20));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(21));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(22));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(23));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(24));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(25));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(26));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(27));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(28));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(29));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(30));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(31));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(32));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(33));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(34));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(35));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(36));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(37));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(38));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(39));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(40));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(41));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(42));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(43));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(44));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(45));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(46));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(47));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(48));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(49));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(50));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(51));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(52));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(53));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(54));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(55));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(56));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(57));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(58));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(59));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(60));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(61));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(62));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(63));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(64));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(65));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(66));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(67));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(68));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(69));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(70));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(71));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(72));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(73));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(74));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(75));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(76));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(77));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(78));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(79));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(80));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(81));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(82));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(83));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(84));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(85));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(86));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(87));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(88));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(89));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(90));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(91));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(92));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(93));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(94));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(95));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(96));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(97));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(98));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(99));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(100));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(101));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(102));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(103));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(104));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(105));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(106));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(107));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(108));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(109));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(110));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(111));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(112));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(113));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(114));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(115));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(116));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(117));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(118));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(119));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(120));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(121));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(122));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(123));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(124));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(125));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(126));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(127));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_char_128(data : std_logic_vector) return char_128 is
        variable rv : char_128;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(16) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(17) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(18) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(19) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(20) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(21) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(22) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(23) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(24) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(25) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(26) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(27) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(28) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(29) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(30) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(31) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(32) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(33) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(34) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(35) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(36) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(37) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(38) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(39) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(40) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(41) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(42) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(43) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(44) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(45) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(46) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(47) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(48) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(49) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(50) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(51) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(52) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(53) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(54) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(55) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(56) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(57) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(58) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(59) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(60) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(61) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(62) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(63) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(64) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(65) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(66) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(67) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(68) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(69) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(70) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(71) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(72) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(73) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(74) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(75) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(76) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(77) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(78) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(79) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(80) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(81) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(82) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(83) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(84) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(85) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(86) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(87) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(88) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(89) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(90) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(91) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(92) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(93) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(94) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(95) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(96) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(97) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(98) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(99) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(100) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(101) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(102) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(103) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(104) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(105) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(106) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(107) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(108) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(109) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(110) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(111) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(112) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(113) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(114) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(115) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(116) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(117) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(118) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(119) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(120) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(121) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(122) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(123) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(124) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(125) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(126) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(127) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function char_2_128_to_slv(data : char_2_128) return std_logic_vector is
        variable rv : std_logic_vector(char_2_128_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+char_128_SLV_LEN)-1 downto pos) := char_128_to_slv(data(0));
            pos := pos + char_128_SLV_LEN;
    
            rv((pos+char_128_SLV_LEN)-1 downto pos) := char_128_to_slv(data(1));
            pos := pos + char_128_SLV_LEN;
    
          return rv;
      end function;
    
      function slv_to_char_2_128(data : std_logic_vector) return char_2_128 is
        variable rv : char_2_128;
        variable elem_slv : std_logic_vector(char_128_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+char_128_SLV_LEN)-1 downto pos);
            rv(0) := slv_to_char_128(elem_slv);
            pos := pos + char_128_SLV_LEN;
    
            elem_slv := data((pos+char_128_SLV_LEN)-1 downto pos);
            rv(1) := slv_to_char_128(elem_slv);
            pos := pos + char_128_SLV_LEN;
    
          return rv;
      end function;
    
      function uint32_t_2_to_slv(data : uint32_t_2) return std_logic_vector is
        variable rv : std_logic_vector(uint32_t_2_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 32;
    
          return rv;
      end function;
    
      function slv_to_uint32_t_2(data : std_logic_vector) return uint32_t_2 is
        variable rv : uint32_t_2;
        variable elem_slv : std_logic_vector(32-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 32;
    
          return rv;
      end function;
    
      function uint8_t_144_to_slv(data : uint8_t_144) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_144_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(16));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(17));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(18));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(19));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(20));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(21));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(22));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(23));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(24));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(25));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(26));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(27));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(28));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(29));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(30));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(31));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(32));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(33));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(34));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(35));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(36));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(37));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(38));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(39));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(40));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(41));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(42));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(43));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(44));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(45));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(46));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(47));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(48));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(49));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(50));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(51));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(52));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(53));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(54));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(55));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(56));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(57));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(58));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(59));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(60));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(61));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(62));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(63));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(64));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(65));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(66));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(67));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(68));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(69));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(70));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(71));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(72));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(73));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(74));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(75));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(76));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(77));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(78));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(79));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(80));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(81));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(82));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(83));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(84));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(85));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(86));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(87));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(88));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(89));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(90));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(91));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(92));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(93));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(94));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(95));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(96));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(97));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(98));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(99));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(100));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(101));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(102));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(103));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(104));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(105));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(106));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(107));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(108));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(109));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(110));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(111));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(112));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(113));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(114));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(115));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(116));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(117));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(118));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(119));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(120));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(121));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(122));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(123));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(124));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(125));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(126));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(127));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(128));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(129));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(130));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(131));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(132));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(133));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(134));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(135));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(136));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(137));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(138));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(139));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(140));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(141));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(142));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(143));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_144(data : std_logic_vector) return uint8_t_144 is
        variable rv : uint8_t_144;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(16) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(17) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(18) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(19) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(20) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(21) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(22) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(23) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(24) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(25) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(26) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(27) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(28) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(29) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(30) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(31) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(32) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(33) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(34) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(35) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(36) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(37) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(38) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(39) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(40) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(41) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(42) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(43) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(44) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(45) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(46) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(47) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(48) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(49) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(50) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(51) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(52) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(53) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(54) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(55) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(56) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(57) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(58) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(59) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(60) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(61) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(62) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(63) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(64) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(65) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(66) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(67) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(68) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(69) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(70) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(71) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(72) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(73) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(74) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(75) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(76) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(77) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(78) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(79) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(80) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(81) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(82) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(83) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(84) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(85) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(86) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(87) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(88) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(89) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(90) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(91) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(92) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(93) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(94) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(95) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(96) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(97) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(98) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(99) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(100) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(101) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(102) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(103) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(104) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(105) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(106) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(107) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(108) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(109) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(110) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(111) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(112) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(113) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(114) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(115) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(116) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(117) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(118) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(119) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(120) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(121) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(122) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(123) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(124) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(125) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(126) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(127) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(128) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(129) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(130) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(131) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(132) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(133) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(134) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(135) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(136) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(137) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(138) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(139) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(140) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(141) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(142) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(143) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function uint8_t_2_144_to_slv(data : uint8_t_2_144) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_2_144_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+uint8_t_144_SLV_LEN)-1 downto pos) := uint8_t_144_to_slv(data(0));
            pos := pos + uint8_t_144_SLV_LEN;
    
            rv((pos+uint8_t_144_SLV_LEN)-1 downto pos) := uint8_t_144_to_slv(data(1));
            pos := pos + uint8_t_144_SLV_LEN;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_2_144(data : std_logic_vector) return uint8_t_2_144 is
        variable rv : uint8_t_2_144;
        variable elem_slv : std_logic_vector(uint8_t_144_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+uint8_t_144_SLV_LEN)-1 downto pos);
            rv(0) := slv_to_uint8_t_144(elem_slv);
            pos := pos + uint8_t_144_SLV_LEN;
    
            elem_slv := data((pos+uint8_t_144_SLV_LEN)-1 downto pos);
            rv(1) := slv_to_uint8_t_144(elem_slv);
            pos := pos + uint8_t_144_SLV_LEN;
    
          return rv;
      end function;
    
      function uint8_t_1_to_slv(data : uint8_t_1) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_1_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_1(data : std_logic_vector) return uint8_t_1 is
        variable rv : uint8_t_1;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function uint1_t_1_to_slv(data : uint1_t_1) return std_logic_vector is
        variable rv : std_logic_vector(uint1_t_1_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 1;
    
          return rv;
      end function;
    
      function slv_to_uint1_t_1(data : std_logic_vector) return uint1_t_1 is
        variable rv : uint1_t_1;
        variable elem_slv : std_logic_vector(1-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 1;
    
          return rv;
      end function;
    
      function uint8_t_2_to_slv(data : uint8_t_2) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_2_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_2(data : std_logic_vector) return uint8_t_2 is
        variable rv : uint8_t_2;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function uint1_t_2_to_slv(data : uint1_t_2) return std_logic_vector is
        variable rv : std_logic_vector(uint1_t_2_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 1;
    
          return rv;
      end function;
    
      function slv_to_uint1_t_2(data : std_logic_vector) return uint1_t_2 is
        variable rv : uint1_t_2;
        variable elem_slv : std_logic_vector(1-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 1;
    
          return rv;
      end function;
    
      function uint8_t_4_to_slv(data : uint8_t_4) return std_logic_vector is
        variable rv : std_logic_vector(uint8_t_4_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 8;
    
            rv((pos+8)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 8;
    
          return rv;
      end function;
    
      function slv_to_uint8_t_4(data : std_logic_vector) return uint8_t_4 is
        variable rv : uint8_t_4;
        variable elem_slv : std_logic_vector(8-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 8;
    
            elem_slv := data((pos+8)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 8;
    
          return rv;
      end function;
    
      function uint1_t_4_to_slv(data : uint1_t_4) return std_logic_vector is
        variable rv : std_logic_vector(uint1_t_4_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 1;
    
          return rv;
      end function;
    
      function slv_to_uint1_t_4(data : std_logic_vector) return uint1_t_4 is
        variable rv : uint1_t_4;
        variable elem_slv : std_logic_vector(1-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 1;
    
          return rv;
      end function;
    
      function uint1_t_8_to_slv(data : uint1_t_8) return std_logic_vector is
        variable rv : std_logic_vector(uint1_t_8_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 1;
    
          return rv;
      end function;
    
      function slv_to_uint1_t_8(data : std_logic_vector) return uint1_t_8 is
        variable rv : uint1_t_8;
        variable elem_slv : std_logic_vector(1-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 1;
    
          return rv;
      end function;
    
      function uint1_t_32_to_slv(data : uint1_t_32) return std_logic_vector is
        variable rv : std_logic_vector(uint1_t_32_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(16));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(17));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(18));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(19));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(20));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(21));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(22));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(23));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(24));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(25));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(26));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(27));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(28));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(29));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(30));
            pos := pos + 1;
    
            rv((pos+1)-1 downto pos) := std_logic_vector(data(31));
            pos := pos + 1;
    
          return rv;
      end function;
    
      function slv_to_uint1_t_32(data : std_logic_vector) return uint1_t_32 is
        variable rv : uint1_t_32;
        variable elem_slv : std_logic_vector(1-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(16) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(17) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(18) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(19) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(20) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(21) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(22) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(23) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(24) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(25) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(26) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(27) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(28) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(29) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(30) := unsigned(elem_slv);
            pos := pos + 1;
    
            elem_slv := data((pos+1)-1 downto pos);
            rv(31) := unsigned(elem_slv);
            pos := pos + 1;
    
          return rv;
      end function;
    
      function uint32_t_16_to_slv(data : uint32_t_16) return std_logic_vector is
        variable rv : std_logic_vector(uint32_t_16_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(0));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(1));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(2));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(3));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(4));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(5));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(6));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(7));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(8));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(9));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(10));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(11));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(12));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(13));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(14));
            pos := pos + 32;
    
            rv((pos+32)-1 downto pos) := std_logic_vector(data(15));
            pos := pos + 32;
    
          return rv;
      end function;
    
      function slv_to_uint32_t_16(data : std_logic_vector) return uint32_t_16 is
        variable rv : uint32_t_16;
        variable elem_slv : std_logic_vector(32-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(0) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(1) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(2) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(3) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(4) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(5) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(6) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(7) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(8) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(9) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(10) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(11) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(12) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(13) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(14) := unsigned(elem_slv);
            pos := pos + 32;
    
            elem_slv := data((pos+32)-1 downto pos);
            rv(15) := unsigned(elem_slv);
            pos := pos + 32;
    
          return rv;
      end function;
    
  function axis8_t_to_slv(data : axis8_t) return std_logic_vector is
    variable rv : std_logic_vector(axis8_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_1_SLV_LEN)-1 downto pos) := uint8_t_1_to_slv(data.tdata);
        pos := pos + uint8_t_1_SLV_LEN;

        rv((pos+uint1_t_1_SLV_LEN)-1 downto pos) := uint1_t_1_to_slv(data.tkeep);
        pos := pos + uint1_t_1_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.tlast);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis8_t(data : std_logic_vector) return axis8_t is
    variable rv : axis8_t;
    variable pos : integer := 0;
    variable tdata_slv : std_logic_vector(uint8_t_1_SLV_LEN-1 downto 0);
    variable tkeep_slv : std_logic_vector(uint1_t_1_SLV_LEN-1 downto 0);
    variable tlast_slv : std_logic_vector(1-1 downto 0);
  begin

        tdata_slv := data((pos+uint8_t_1_SLV_LEN)-1 downto pos);
        rv.tdata := slv_to_uint8_t_1(tdata_slv);
        pos := pos + uint8_t_1_SLV_LEN;

        tkeep_slv := data((pos+uint1_t_1_SLV_LEN)-1 downto pos);
        rv.tkeep := slv_to_uint1_t_1(tkeep_slv);
        pos := pos + uint1_t_1_SLV_LEN;

        tlast_slv := data((pos+1)-1 downto pos);
        rv.tlast := unsigned(tlast_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis8_t_stream_t_to_slv(data : axis8_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(axis8_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis8_t_SLV_LEN)-1 downto pos) := axis8_t_to_slv(data.data);
        pos := pos + axis8_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis8_t_stream_t(data : std_logic_vector) return axis8_t_stream_t is
    variable rv : axis8_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(axis8_t_SLV_LEN-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+axis8_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_axis8_t(data_slv);
        pos := pos + axis8_t_SLV_LEN;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis16_t_to_slv(data : axis16_t) return std_logic_vector is
    variable rv : std_logic_vector(axis16_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_2_SLV_LEN)-1 downto pos) := uint8_t_2_to_slv(data.tdata);
        pos := pos + uint8_t_2_SLV_LEN;

        rv((pos+uint1_t_2_SLV_LEN)-1 downto pos) := uint1_t_2_to_slv(data.tkeep);
        pos := pos + uint1_t_2_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.tlast);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis16_t(data : std_logic_vector) return axis16_t is
    variable rv : axis16_t;
    variable pos : integer := 0;
    variable tdata_slv : std_logic_vector(uint8_t_2_SLV_LEN-1 downto 0);
    variable tkeep_slv : std_logic_vector(uint1_t_2_SLV_LEN-1 downto 0);
    variable tlast_slv : std_logic_vector(1-1 downto 0);
  begin

        tdata_slv := data((pos+uint8_t_2_SLV_LEN)-1 downto pos);
        rv.tdata := slv_to_uint8_t_2(tdata_slv);
        pos := pos + uint8_t_2_SLV_LEN;

        tkeep_slv := data((pos+uint1_t_2_SLV_LEN)-1 downto pos);
        rv.tkeep := slv_to_uint1_t_2(tkeep_slv);
        pos := pos + uint1_t_2_SLV_LEN;

        tlast_slv := data((pos+1)-1 downto pos);
        rv.tlast := unsigned(tlast_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis16_t_stream_t_to_slv(data : axis16_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(axis16_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis16_t_SLV_LEN)-1 downto pos) := axis16_t_to_slv(data.data);
        pos := pos + axis16_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis16_t_stream_t(data : std_logic_vector) return axis16_t_stream_t is
    variable rv : axis16_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(axis16_t_SLV_LEN-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+axis16_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_axis16_t(data_slv);
        pos := pos + axis16_t_SLV_LEN;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis32_t_to_slv(data : axis32_t) return std_logic_vector is
    variable rv : std_logic_vector(axis32_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_4_SLV_LEN)-1 downto pos) := uint8_t_4_to_slv(data.tdata);
        pos := pos + uint8_t_4_SLV_LEN;

        rv((pos+uint1_t_4_SLV_LEN)-1 downto pos) := uint1_t_4_to_slv(data.tkeep);
        pos := pos + uint1_t_4_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.tlast);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis32_t(data : std_logic_vector) return axis32_t is
    variable rv : axis32_t;
    variable pos : integer := 0;
    variable tdata_slv : std_logic_vector(uint8_t_4_SLV_LEN-1 downto 0);
    variable tkeep_slv : std_logic_vector(uint1_t_4_SLV_LEN-1 downto 0);
    variable tlast_slv : std_logic_vector(1-1 downto 0);
  begin

        tdata_slv := data((pos+uint8_t_4_SLV_LEN)-1 downto pos);
        rv.tdata := slv_to_uint8_t_4(tdata_slv);
        pos := pos + uint8_t_4_SLV_LEN;

        tkeep_slv := data((pos+uint1_t_4_SLV_LEN)-1 downto pos);
        rv.tkeep := slv_to_uint1_t_4(tkeep_slv);
        pos := pos + uint1_t_4_SLV_LEN;

        tlast_slv := data((pos+1)-1 downto pos);
        rv.tlast := unsigned(tlast_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis32_t_stream_t_to_slv(data : axis32_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(axis32_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis32_t_SLV_LEN)-1 downto pos) := axis32_t_to_slv(data.data);
        pos := pos + axis32_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis32_t_stream_t(data : std_logic_vector) return axis32_t_stream_t is
    variable rv : axis32_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(axis32_t_SLV_LEN-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+axis32_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_axis32_t(data_slv);
        pos := pos + axis32_t_SLV_LEN;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis64_t_to_slv(data : axis64_t) return std_logic_vector is
    variable rv : std_logic_vector(axis64_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_8_SLV_LEN)-1 downto pos) := uint8_t_8_to_slv(data.tdata);
        pos := pos + uint8_t_8_SLV_LEN;

        rv((pos+uint1_t_8_SLV_LEN)-1 downto pos) := uint1_t_8_to_slv(data.tkeep);
        pos := pos + uint1_t_8_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.tlast);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis64_t(data : std_logic_vector) return axis64_t is
    variable rv : axis64_t;
    variable pos : integer := 0;
    variable tdata_slv : std_logic_vector(uint8_t_8_SLV_LEN-1 downto 0);
    variable tkeep_slv : std_logic_vector(uint1_t_8_SLV_LEN-1 downto 0);
    variable tlast_slv : std_logic_vector(1-1 downto 0);
  begin

        tdata_slv := data((pos+uint8_t_8_SLV_LEN)-1 downto pos);
        rv.tdata := slv_to_uint8_t_8(tdata_slv);
        pos := pos + uint8_t_8_SLV_LEN;

        tkeep_slv := data((pos+uint1_t_8_SLV_LEN)-1 downto pos);
        rv.tkeep := slv_to_uint1_t_8(tkeep_slv);
        pos := pos + uint1_t_8_SLV_LEN;

        tlast_slv := data((pos+1)-1 downto pos);
        rv.tlast := unsigned(tlast_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis64_t_stream_t_to_slv(data : axis64_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(axis64_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis64_t_SLV_LEN)-1 downto pos) := axis64_t_to_slv(data.data);
        pos := pos + axis64_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis64_t_stream_t(data : std_logic_vector) return axis64_t_stream_t is
    variable rv : axis64_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(axis64_t_SLV_LEN-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+axis64_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_axis64_t(data_slv);
        pos := pos + axis64_t_SLV_LEN;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis128_t_to_slv(data : axis128_t) return std_logic_vector is
    variable rv : std_logic_vector(axis128_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_16_SLV_LEN)-1 downto pos) := uint8_t_16_to_slv(data.tdata);
        pos := pos + uint8_t_16_SLV_LEN;

        rv((pos+uint1_t_16_SLV_LEN)-1 downto pos) := uint1_t_16_to_slv(data.tkeep);
        pos := pos + uint1_t_16_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.tlast);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis128_t(data : std_logic_vector) return axis128_t is
    variable rv : axis128_t;
    variable pos : integer := 0;
    variable tdata_slv : std_logic_vector(uint8_t_16_SLV_LEN-1 downto 0);
    variable tkeep_slv : std_logic_vector(uint1_t_16_SLV_LEN-1 downto 0);
    variable tlast_slv : std_logic_vector(1-1 downto 0);
  begin

        tdata_slv := data((pos+uint8_t_16_SLV_LEN)-1 downto pos);
        rv.tdata := slv_to_uint8_t_16(tdata_slv);
        pos := pos + uint8_t_16_SLV_LEN;

        tkeep_slv := data((pos+uint1_t_16_SLV_LEN)-1 downto pos);
        rv.tkeep := slv_to_uint1_t_16(tkeep_slv);
        pos := pos + uint1_t_16_SLV_LEN;

        tlast_slv := data((pos+1)-1 downto pos);
        rv.tlast := unsigned(tlast_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis128_t_stream_t_to_slv(data : axis128_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(axis128_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis128_t_SLV_LEN)-1 downto pos) := axis128_t_to_slv(data.data);
        pos := pos + axis128_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis128_t_stream_t(data : std_logic_vector) return axis128_t_stream_t is
    variable rv : axis128_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(axis128_t_SLV_LEN-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+axis128_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_axis128_t(data_slv);
        pos := pos + axis128_t_SLV_LEN;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis256_t_to_slv(data : axis256_t) return std_logic_vector is
    variable rv : std_logic_vector(axis256_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_32_SLV_LEN)-1 downto pos) := uint8_t_32_to_slv(data.tdata);
        pos := pos + uint8_t_32_SLV_LEN;

        rv((pos+uint1_t_32_SLV_LEN)-1 downto pos) := uint1_t_32_to_slv(data.tkeep);
        pos := pos + uint1_t_32_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.tlast);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis256_t(data : std_logic_vector) return axis256_t is
    variable rv : axis256_t;
    variable pos : integer := 0;
    variable tdata_slv : std_logic_vector(uint8_t_32_SLV_LEN-1 downto 0);
    variable tkeep_slv : std_logic_vector(uint1_t_32_SLV_LEN-1 downto 0);
    variable tlast_slv : std_logic_vector(1-1 downto 0);
  begin

        tdata_slv := data((pos+uint8_t_32_SLV_LEN)-1 downto pos);
        rv.tdata := slv_to_uint8_t_32(tdata_slv);
        pos := pos + uint8_t_32_SLV_LEN;

        tkeep_slv := data((pos+uint1_t_32_SLV_LEN)-1 downto pos);
        rv.tkeep := slv_to_uint1_t_32(tkeep_slv);
        pos := pos + uint1_t_32_SLV_LEN;

        tlast_slv := data((pos+1)-1 downto pos);
        rv.tlast := unsigned(tlast_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis256_t_stream_t_to_slv(data : axis256_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(axis256_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis256_t_SLV_LEN)-1 downto pos) := axis256_t_to_slv(data.data);
        pos := pos + axis256_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis256_t_stream_t(data : std_logic_vector) return axis256_t_stream_t is
    variable rv : axis256_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(axis256_t_SLV_LEN-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+axis256_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_axis256_t(data_slv);
        pos := pos + axis256_t_SLV_LEN;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis512_t_to_slv(data : axis512_t) return std_logic_vector is
    variable rv : std_logic_vector(axis512_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_64_SLV_LEN)-1 downto pos) := uint8_t_64_to_slv(data.tdata);
        pos := pos + uint8_t_64_SLV_LEN;

        rv((pos+uint1_t_64_SLV_LEN)-1 downto pos) := uint1_t_64_to_slv(data.tkeep);
        pos := pos + uint1_t_64_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.tlast);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis512_t(data : std_logic_vector) return axis512_t is
    variable rv : axis512_t;
    variable pos : integer := 0;
    variable tdata_slv : std_logic_vector(uint8_t_64_SLV_LEN-1 downto 0);
    variable tkeep_slv : std_logic_vector(uint1_t_64_SLV_LEN-1 downto 0);
    variable tlast_slv : std_logic_vector(1-1 downto 0);
  begin

        tdata_slv := data((pos+uint8_t_64_SLV_LEN)-1 downto pos);
        rv.tdata := slv_to_uint8_t_64(tdata_slv);
        pos := pos + uint8_t_64_SLV_LEN;

        tkeep_slv := data((pos+uint1_t_64_SLV_LEN)-1 downto pos);
        rv.tkeep := slv_to_uint1_t_64(tkeep_slv);
        pos := pos + uint1_t_64_SLV_LEN;

        tlast_slv := data((pos+1)-1 downto pos);
        rv.tlast := unsigned(tlast_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis512_t_stream_t_to_slv(data : axis512_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(axis512_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis512_t_SLV_LEN)-1 downto pos) := axis512_t_to_slv(data.data);
        pos := pos + axis512_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis512_t_stream_t(data : std_logic_vector) return axis512_t_stream_t is
    variable rv : axis512_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(axis512_t_SLV_LEN-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+axis512_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_axis512_t(data_slv);
        pos := pos + axis512_t_SLV_LEN;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis8_to_axis32_t_to_slv(data : axis8_to_axis32_t) return std_logic_vector is
    variable rv : std_logic_vector(axis8_to_axis32_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis32_t_stream_t_SLV_LEN)-1 downto pos) := axis32_t_stream_t_to_slv(data.axis_out);
        pos := pos + axis32_t_stream_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.axis_in_ready);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis8_to_axis32_t(data : std_logic_vector) return axis8_to_axis32_t is
    variable rv : axis8_to_axis32_t;
    variable pos : integer := 0;
    variable axis_out_slv : std_logic_vector(axis32_t_stream_t_SLV_LEN-1 downto 0);
    variable axis_in_ready_slv : std_logic_vector(1-1 downto 0);
  begin

        axis_out_slv := data((pos+axis32_t_stream_t_SLV_LEN)-1 downto pos);
        rv.axis_out := slv_to_axis32_t_stream_t(axis_out_slv);
        pos := pos + axis32_t_stream_t_SLV_LEN;

        axis_in_ready_slv := data((pos+1)-1 downto pos);
        rv.axis_in_ready := unsigned(axis_in_ready_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis32_to_axis8_t_to_slv(data : axis32_to_axis8_t) return std_logic_vector is
    variable rv : std_logic_vector(axis32_to_axis8_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis8_t_stream_t_SLV_LEN)-1 downto pos) := axis8_t_stream_t_to_slv(data.axis_out);
        pos := pos + axis8_t_stream_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.axis_in_ready);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis32_to_axis8_t(data : std_logic_vector) return axis32_to_axis8_t is
    variable rv : axis32_to_axis8_t;
    variable pos : integer := 0;
    variable axis_out_slv : std_logic_vector(axis8_t_stream_t_SLV_LEN-1 downto 0);
    variable axis_in_ready_slv : std_logic_vector(1-1 downto 0);
  begin

        axis_out_slv := data((pos+axis8_t_stream_t_SLV_LEN)-1 downto pos);
        rv.axis_out := slv_to_axis8_t_stream_t(axis_out_slv);
        pos := pos + axis8_t_stream_t_SLV_LEN;

        axis_in_ready_slv := data((pos+1)-1 downto pos);
        rv.axis_in_ready := unsigned(axis_in_ready_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis128_to_axis512_t_to_slv(data : axis128_to_axis512_t) return std_logic_vector is
    variable rv : std_logic_vector(axis128_to_axis512_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis512_t_stream_t_SLV_LEN)-1 downto pos) := axis512_t_stream_t_to_slv(data.axis_out);
        pos := pos + axis512_t_stream_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.axis_in_ready);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis128_to_axis512_t(data : std_logic_vector) return axis128_to_axis512_t is
    variable rv : axis128_to_axis512_t;
    variable pos : integer := 0;
    variable axis_out_slv : std_logic_vector(axis512_t_stream_t_SLV_LEN-1 downto 0);
    variable axis_in_ready_slv : std_logic_vector(1-1 downto 0);
  begin

        axis_out_slv := data((pos+axis512_t_stream_t_SLV_LEN)-1 downto pos);
        rv.axis_out := slv_to_axis512_t_stream_t(axis_out_slv);
        pos := pos + axis512_t_stream_t_SLV_LEN;

        axis_in_ready_slv := data((pos+1)-1 downto pos);
        rv.axis_in_ready := unsigned(axis_in_ready_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis512_to_axis128_t_to_slv(data : axis512_to_axis128_t) return std_logic_vector is
    variable rv : std_logic_vector(axis512_to_axis128_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos) := axis128_t_stream_t_to_slv(data.axis_out);
        pos := pos + axis128_t_stream_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.axis_in_ready);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis512_to_axis128_t(data : std_logic_vector) return axis512_to_axis128_t is
    variable rv : axis512_to_axis128_t;
    variable pos : integer := 0;
    variable axis_out_slv : std_logic_vector(axis128_t_stream_t_SLV_LEN-1 downto 0);
    variable axis_in_ready_slv : std_logic_vector(1-1 downto 0);
  begin

        axis_out_slv := data((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos);
        rv.axis_out := slv_to_axis128_t_stream_t(axis_out_slv);
        pos := pos + axis128_t_stream_t_SLV_LEN;

        axis_in_ready_slv := data((pos+1)-1 downto pos);
        rv.axis_in_ready := unsigned(axis_in_ready_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis8_max_len_limiter_t_to_slv(data : axis8_max_len_limiter_t) return std_logic_vector is
    variable rv : std_logic_vector(axis8_max_len_limiter_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis8_t_stream_t_SLV_LEN)-1 downto pos) := axis8_t_stream_t_to_slv(data.out_stream);
        pos := pos + axis8_t_stream_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.ready_for_in_stream);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis8_max_len_limiter_t(data : std_logic_vector) return axis8_max_len_limiter_t is
    variable rv : axis8_max_len_limiter_t;
    variable pos : integer := 0;
    variable out_stream_slv : std_logic_vector(axis8_t_stream_t_SLV_LEN-1 downto 0);
    variable ready_for_in_stream_slv : std_logic_vector(1-1 downto 0);
  begin

        out_stream_slv := data((pos+axis8_t_stream_t_SLV_LEN)-1 downto pos);
        rv.out_stream := slv_to_axis8_t_stream_t(out_stream_slv);
        pos := pos + axis8_t_stream_t_SLV_LEN;

        ready_for_in_stream_slv := data((pos+1)-1 downto pos);
        rv.ready_for_in_stream := unsigned(ready_for_in_stream_slv);
        pos := pos + 1;

      return rv;
  end function;

  function axis32_max_len_limiter_t_to_slv(data : axis32_max_len_limiter_t) return std_logic_vector is
    variable rv : std_logic_vector(axis32_max_len_limiter_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis32_t_stream_t_SLV_LEN)-1 downto pos) := axis32_t_stream_t_to_slv(data.out_stream);
        pos := pos + axis32_t_stream_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.ready_for_in_stream);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_axis32_max_len_limiter_t(data : std_logic_vector) return axis32_max_len_limiter_t is
    variable rv : axis32_max_len_limiter_t;
    variable pos : integer := 0;
    variable out_stream_slv : std_logic_vector(axis32_t_stream_t_SLV_LEN-1 downto 0);
    variable ready_for_in_stream_slv : std_logic_vector(1-1 downto 0);
  begin

        out_stream_slv := data((pos+axis32_t_stream_t_SLV_LEN)-1 downto pos);
        rv.out_stream := slv_to_axis32_t_stream_t(out_stream_slv);
        pos := pos + axis32_t_stream_t_SLV_LEN;

        ready_for_in_stream_slv := data((pos+1)-1 downto pos);
        rv.ready_for_in_stream := unsigned(ready_for_in_stream_slv);
        pos := pos + 1;

      return rv;
  end function;

  function chacha20_state_to_slv(data : chacha20_state) return std_logic_vector is
    variable rv : std_logic_vector(chacha20_state_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint32_t_16_SLV_LEN)-1 downto pos) := uint32_t_16_to_slv(data.state);
        pos := pos + uint32_t_16_SLV_LEN;

      return rv;
  end function;

  function slv_to_chacha20_state(data : std_logic_vector) return chacha20_state is
    variable rv : chacha20_state;
    variable pos : integer := 0;
    variable state_slv : std_logic_vector(uint32_t_16_SLV_LEN-1 downto 0);
  begin

        state_slv := data((pos+uint32_t_16_SLV_LEN)-1 downto pos);
        rv.state := slv_to_uint32_t_16(state_slv);
        pos := pos + uint32_t_16_SLV_LEN;

      return rv;
  end function;

  function chacha20_decrypt_loop_body_in_t_to_slv(data : chacha20_decrypt_loop_body_in_t) return std_logic_vector is
    variable rv : std_logic_vector(chacha20_decrypt_loop_body_in_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis512_t_SLV_LEN)-1 downto pos) := axis512_t_to_slv(data.axis_in);
        pos := pos + axis512_t_SLV_LEN;

        rv((pos+uint8_t_32_SLV_LEN)-1 downto pos) := uint8_t_32_to_slv(data.key);
        pos := pos + uint8_t_32_SLV_LEN;

        rv((pos+uint8_t_12_SLV_LEN)-1 downto pos) := uint8_t_12_to_slv(data.nonce);
        pos := pos + uint8_t_12_SLV_LEN;

        rv((pos+32)-1 downto pos) := std_logic_vector(data.counter);
        pos := pos + 32;

      return rv;
  end function;

  function slv_to_chacha20_decrypt_loop_body_in_t(data : std_logic_vector) return chacha20_decrypt_loop_body_in_t is
    variable rv : chacha20_decrypt_loop_body_in_t;
    variable pos : integer := 0;
    variable axis_in_slv : std_logic_vector(axis512_t_SLV_LEN-1 downto 0);
    variable key_slv : std_logic_vector(uint8_t_32_SLV_LEN-1 downto 0);
    variable nonce_slv : std_logic_vector(uint8_t_12_SLV_LEN-1 downto 0);
    variable counter_slv : std_logic_vector(32-1 downto 0);
  begin

        axis_in_slv := data((pos+axis512_t_SLV_LEN)-1 downto pos);
        rv.axis_in := slv_to_axis512_t(axis_in_slv);
        pos := pos + axis512_t_SLV_LEN;

        key_slv := data((pos+uint8_t_32_SLV_LEN)-1 downto pos);
        rv.key := slv_to_uint8_t_32(key_slv);
        pos := pos + uint8_t_32_SLV_LEN;

        nonce_slv := data((pos+uint8_t_12_SLV_LEN)-1 downto pos);
        rv.nonce := slv_to_uint8_t_12(nonce_slv);
        pos := pos + uint8_t_12_SLV_LEN;

        counter_slv := data((pos+32)-1 downto pos);
        rv.counter := unsigned(counter_slv);
        pos := pos + 32;

      return rv;
  end function;

  function chacha20_decrypt_loop_body_in_t_stream_t_to_slv(data : chacha20_decrypt_loop_body_in_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(chacha20_decrypt_loop_body_in_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+chacha20_decrypt_loop_body_in_t_SLV_LEN)-1 downto pos) := chacha20_decrypt_loop_body_in_t_to_slv(data.data);
        pos := pos + chacha20_decrypt_loop_body_in_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_chacha20_decrypt_loop_body_in_t_stream_t(data : std_logic_vector) return chacha20_decrypt_loop_body_in_t_stream_t is
    variable rv : chacha20_decrypt_loop_body_in_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(chacha20_decrypt_loop_body_in_t_SLV_LEN-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+chacha20_decrypt_loop_body_in_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_chacha20_decrypt_loop_body_in_t(data_slv);
        pos := pos + chacha20_decrypt_loop_body_in_t_SLV_LEN;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function uint256_t_stream_t_to_slv(data : uint256_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(uint256_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+256)-1 downto pos) := std_logic_vector(data.data);
        pos := pos + 256;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_uint256_t_stream_t(data : std_logic_vector) return uint256_t_stream_t is
    variable rv : uint256_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(256-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+256)-1 downto pos);
        rv.data := unsigned(data_slv);
        pos := pos + 256;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function uint128_t_stream_t_to_slv(data : uint128_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(uint128_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+128)-1 downto pos) := std_logic_vector(data.data);
        pos := pos + 128;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_uint128_t_stream_t(data : std_logic_vector) return uint128_t_stream_t is
    variable rv : uint128_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(128-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+128)-1 downto pos);
        rv.data := unsigned(data_slv);
        pos := pos + 128;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function u320_t_to_slv(data : u320_t) return std_logic_vector is
    variable rv : std_logic_vector(u320_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint64_t_5_SLV_LEN)-1 downto pos) := uint64_t_5_to_slv(data.limbs);
        pos := pos + uint64_t_5_SLV_LEN;

      return rv;
  end function;

  function slv_to_u320_t(data : std_logic_vector) return u320_t is
    variable rv : u320_t;
    variable pos : integer := 0;
    variable limbs_slv : std_logic_vector(uint64_t_5_SLV_LEN-1 downto 0);
  begin

        limbs_slv := data((pos+uint64_t_5_SLV_LEN)-1 downto pos);
        rv.limbs := slv_to_uint64_t_5(limbs_slv);
        pos := pos + uint64_t_5_SLV_LEN;

      return rv;
  end function;

  function u8_16_t_to_slv(data : u8_16_t) return std_logic_vector is
    variable rv : std_logic_vector(u8_16_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_16_SLV_LEN)-1 downto pos) := uint8_t_16_to_slv(data.bytes);
        pos := pos + uint8_t_16_SLV_LEN;

      return rv;
  end function;

  function slv_to_u8_16_t(data : std_logic_vector) return u8_16_t is
    variable rv : u8_16_t;
    variable pos : integer := 0;
    variable bytes_slv : std_logic_vector(uint8_t_16_SLV_LEN-1 downto 0);
  begin

        bytes_slv := data((pos+uint8_t_16_SLV_LEN)-1 downto pos);
        rv.bytes := slv_to_uint8_t_16(bytes_slv);
        pos := pos + uint8_t_16_SLV_LEN;

      return rv;
  end function;

  function poly1305_mac_loop_body_in_t_to_slv(data : poly1305_mac_loop_body_in_t) return std_logic_vector is
    variable rv : std_logic_vector(poly1305_mac_loop_body_in_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_16_SLV_LEN)-1 downto pos) := uint8_t_16_to_slv(data.block_bytes);
        pos := pos + uint8_t_16_SLV_LEN;

        rv((pos+u320_t_SLV_LEN)-1 downto pos) := u320_t_to_slv(data.r);
        pos := pos + u320_t_SLV_LEN;

        rv((pos+u320_t_SLV_LEN)-1 downto pos) := u320_t_to_slv(data.a);
        pos := pos + u320_t_SLV_LEN;

      return rv;
  end function;

  function slv_to_poly1305_mac_loop_body_in_t(data : std_logic_vector) return poly1305_mac_loop_body_in_t is
    variable rv : poly1305_mac_loop_body_in_t;
    variable pos : integer := 0;
    variable block_bytes_slv : std_logic_vector(uint8_t_16_SLV_LEN-1 downto 0);
    variable r_slv : std_logic_vector(u320_t_SLV_LEN-1 downto 0);
    variable a_slv : std_logic_vector(u320_t_SLV_LEN-1 downto 0);
  begin

        block_bytes_slv := data((pos+uint8_t_16_SLV_LEN)-1 downto pos);
        rv.block_bytes := slv_to_uint8_t_16(block_bytes_slv);
        pos := pos + uint8_t_16_SLV_LEN;

        r_slv := data((pos+u320_t_SLV_LEN)-1 downto pos);
        rv.r := slv_to_u320_t(r_slv);
        pos := pos + u320_t_SLV_LEN;

        a_slv := data((pos+u320_t_SLV_LEN)-1 downto pos);
        rv.a := slv_to_u320_t(a_slv);
        pos := pos + u320_t_SLV_LEN;

      return rv;
  end function;

  function chacha20_decrypt_pipeline_no_handshake_in_reg_t_to_slv(data : chacha20_decrypt_pipeline_no_handshake_in_reg_t) return std_logic_vector is
    variable rv : std_logic_vector(chacha20_decrypt_pipeline_no_handshake_in_reg_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+chacha20_decrypt_loop_body_in_t_SLV_LEN)-1 downto pos) := chacha20_decrypt_loop_body_in_t_to_slv(data.data);
        pos := pos + chacha20_decrypt_loop_body_in_t_SLV_LEN;

        rv((pos+8)-1 downto pos) := std_logic_vector(data.id);
        pos := pos + 8;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_chacha20_decrypt_pipeline_no_handshake_in_reg_t(data : std_logic_vector) return chacha20_decrypt_pipeline_no_handshake_in_reg_t is
    variable rv : chacha20_decrypt_pipeline_no_handshake_in_reg_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(chacha20_decrypt_loop_body_in_t_SLV_LEN-1 downto 0);
    variable id_slv : std_logic_vector(8-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+chacha20_decrypt_loop_body_in_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_chacha20_decrypt_loop_body_in_t(data_slv);
        pos := pos + chacha20_decrypt_loop_body_in_t_SLV_LEN;

        id_slv := data((pos+8)-1 downto pos);
        rv.id := unsigned(id_slv);
        pos := pos + 8;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function chacha20_decrypt_pipeline_no_handshake_out_reg_t_to_slv(data : chacha20_decrypt_pipeline_no_handshake_out_reg_t) return std_logic_vector is
    variable rv : std_logic_vector(chacha20_decrypt_pipeline_no_handshake_out_reg_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis512_t_SLV_LEN)-1 downto pos) := axis512_t_to_slv(data.data);
        pos := pos + axis512_t_SLV_LEN;

        rv((pos+8)-1 downto pos) := std_logic_vector(data.id);
        pos := pos + 8;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_chacha20_decrypt_pipeline_no_handshake_out_reg_t(data : std_logic_vector) return chacha20_decrypt_pipeline_no_handshake_out_reg_t is
    variable rv : chacha20_decrypt_pipeline_no_handshake_out_reg_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(axis512_t_SLV_LEN-1 downto 0);
    variable id_slv : std_logic_vector(8-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+axis512_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_axis512_t(data_slv);
        pos := pos + axis512_t_SLV_LEN;

        id_slv := data((pos+8)-1 downto pos);
        rv.id := unsigned(id_slv);
        pos := pos + 8;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function chacha20_decrypt_pipeline_FIFO_t_to_slv(data : chacha20_decrypt_pipeline_FIFO_t) return std_logic_vector is
    variable rv : std_logic_vector(chacha20_decrypt_pipeline_FIFO_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis512_t_SLV_LEN)-1 downto pos) := axis512_t_to_slv(data.data_out);
        pos := pos + axis512_t_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.data_out_valid);
        pos := pos + 1;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.data_in_ready);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_chacha20_decrypt_pipeline_FIFO_t(data : std_logic_vector) return chacha20_decrypt_pipeline_FIFO_t is
    variable rv : chacha20_decrypt_pipeline_FIFO_t;
    variable pos : integer := 0;
    variable data_out_slv : std_logic_vector(axis512_t_SLV_LEN-1 downto 0);
    variable data_out_valid_slv : std_logic_vector(1-1 downto 0);
    variable data_in_ready_slv : std_logic_vector(1-1 downto 0);
  begin

        data_out_slv := data((pos+axis512_t_SLV_LEN)-1 downto pos);
        rv.data_out := slv_to_axis512_t(data_out_slv);
        pos := pos + axis512_t_SLV_LEN;

        data_out_valid_slv := data((pos+1)-1 downto pos);
        rv.data_out_valid := unsigned(data_out_valid_slv);
        pos := pos + 1;

        data_in_ready_slv := data((pos+1)-1 downto pos);
        rv.data_in_ready := unsigned(data_in_ready_slv);
        pos := pos + 1;

      return rv;
  end function;

  function poly1305_pipeline_in_reg_t_to_slv(data : poly1305_pipeline_in_reg_t) return std_logic_vector is
    variable rv : std_logic_vector(poly1305_pipeline_in_reg_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+poly1305_mac_loop_body_in_t_SLV_LEN)-1 downto pos) := poly1305_mac_loop_body_in_t_to_slv(data.data);
        pos := pos + poly1305_mac_loop_body_in_t_SLV_LEN;

        rv((pos+8)-1 downto pos) := std_logic_vector(data.id);
        pos := pos + 8;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_poly1305_pipeline_in_reg_t(data : std_logic_vector) return poly1305_pipeline_in_reg_t is
    variable rv : poly1305_pipeline_in_reg_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(poly1305_mac_loop_body_in_t_SLV_LEN-1 downto 0);
    variable id_slv : std_logic_vector(8-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+poly1305_mac_loop_body_in_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_poly1305_mac_loop_body_in_t(data_slv);
        pos := pos + poly1305_mac_loop_body_in_t_SLV_LEN;

        id_slv := data((pos+8)-1 downto pos);
        rv.id := unsigned(id_slv);
        pos := pos + 8;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function poly1305_pipeline_out_reg_t_to_slv(data : poly1305_pipeline_out_reg_t) return std_logic_vector is
    variable rv : std_logic_vector(poly1305_pipeline_out_reg_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+u320_t_SLV_LEN)-1 downto pos) := u320_t_to_slv(data.data);
        pos := pos + u320_t_SLV_LEN;

        rv((pos+8)-1 downto pos) := std_logic_vector(data.id);
        pos := pos + 8;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_poly1305_pipeline_out_reg_t(data : std_logic_vector) return poly1305_pipeline_out_reg_t is
    variable rv : poly1305_pipeline_out_reg_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(u320_t_SLV_LEN-1 downto 0);
    variable id_slv : std_logic_vector(8-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+u320_t_SLV_LEN)-1 downto pos);
        rv.data := slv_to_u320_t(data_slv);
        pos := pos + u320_t_SLV_LEN;

        id_slv := data((pos+8)-1 downto pos);
        rv.id := unsigned(id_slv);
        pos := pos + 8;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function uint1_t_stream_t_to_slv(data : uint1_t_stream_t) return std_logic_vector is
    variable rv : std_logic_vector(uint1_t_stream_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+1)-1 downto pos) := std_logic_vector(data.data);
        pos := pos + 1;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_uint1_t_stream_t(data : std_logic_vector) return uint1_t_stream_t is
    variable rv : uint1_t_stream_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(1-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+1)-1 downto pos);
        rv.data := unsigned(data_slv);
        pos := pos + 1;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;

  function verify_fifo_FIFO_write_t_to_slv(data : verify_fifo_FIFO_write_t) return std_logic_vector is
    variable rv : std_logic_vector(verify_fifo_FIFO_write_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+1)-1 downto pos) := std_logic_vector(data.ready);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_verify_fifo_FIFO_write_t(data : std_logic_vector) return verify_fifo_FIFO_write_t is
    variable rv : verify_fifo_FIFO_write_t;
    variable pos : integer := 0;
    variable ready_slv : std_logic_vector(1-1 downto 0);
  begin

        ready_slv := data((pos+1)-1 downto pos);
        rv.ready := unsigned(ready_slv);
        pos := pos + 1;

      return rv;
  end function;

  function uint8_t_array_64_t_to_slv(data : uint8_t_array_64_t) return std_logic_vector is
    variable rv : std_logic_vector(uint8_t_array_64_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_64_SLV_LEN)-1 downto pos) := uint8_t_64_to_slv(data.data);
        pos := pos + uint8_t_64_SLV_LEN;

      return rv;
  end function;

  function slv_to_uint8_t_array_64_t(data : std_logic_vector) return uint8_t_array_64_t is
    variable rv : uint8_t_array_64_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(uint8_t_64_SLV_LEN-1 downto 0);
  begin

        data_slv := data((pos+uint8_t_64_SLV_LEN)-1 downto pos);
        rv.data := slv_to_uint8_t_64(data_slv);
        pos := pos + uint8_t_64_SLV_LEN;

      return rv;
  end function;

  function uint8_t_array_40_t_to_slv(data : uint8_t_array_40_t) return std_logic_vector is
    variable rv : std_logic_vector(uint8_t_array_40_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_40_SLV_LEN)-1 downto pos) := uint8_t_40_to_slv(data.data);
        pos := pos + uint8_t_40_SLV_LEN;

      return rv;
  end function;

  function slv_to_uint8_t_array_40_t(data : std_logic_vector) return uint8_t_array_40_t is
    variable rv : uint8_t_array_40_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(uint8_t_40_SLV_LEN-1 downto 0);
  begin

        data_slv := data((pos+uint8_t_40_SLV_LEN)-1 downto pos);
        rv.data := slv_to_uint8_t_40(data_slv);
        pos := pos + uint8_t_40_SLV_LEN;

      return rv;
  end function;

  function uint8_t_array_8_t_to_slv(data : uint8_t_array_8_t) return std_logic_vector is
    variable rv : std_logic_vector(uint8_t_array_8_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_8_SLV_LEN)-1 downto pos) := uint8_t_8_to_slv(data.data);
        pos := pos + uint8_t_8_SLV_LEN;

      return rv;
  end function;

  function slv_to_uint8_t_array_8_t(data : std_logic_vector) return uint8_t_array_8_t is
    variable rv : uint8_t_array_8_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(uint8_t_8_SLV_LEN-1 downto 0);
  begin

        data_slv := data((pos+uint8_t_8_SLV_LEN)-1 downto pos);
        rv.data := slv_to_uint8_t_8(data_slv);
        pos := pos + uint8_t_8_SLV_LEN;

      return rv;
  end function;

  function uint8_t_array_4_t_to_slv(data : uint8_t_array_4_t) return std_logic_vector is
    variable rv : std_logic_vector(uint8_t_array_4_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_4_SLV_LEN)-1 downto pos) := uint8_t_4_to_slv(data.data);
        pos := pos + uint8_t_4_SLV_LEN;

      return rv;
  end function;

  function slv_to_uint8_t_array_4_t(data : std_logic_vector) return uint8_t_array_4_t is
    variable rv : uint8_t_array_4_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(uint8_t_4_SLV_LEN-1 downto 0);
  begin

        data_slv := data((pos+uint8_t_4_SLV_LEN)-1 downto pos);
        rv.data := slv_to_uint8_t_4(data_slv);
        pos := pos + uint8_t_4_SLV_LEN;

      return rv;
  end function;

  function uint32_t_array_16_t_to_slv(data : uint32_t_array_16_t) return std_logic_vector is
    variable rv : std_logic_vector(uint32_t_array_16_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint32_t_16_SLV_LEN)-1 downto pos) := uint32_t_16_to_slv(data.data);
        pos := pos + uint32_t_16_SLV_LEN;

      return rv;
  end function;

  function slv_to_uint32_t_array_16_t(data : std_logic_vector) return uint32_t_array_16_t is
    variable rv : uint32_t_array_16_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(uint32_t_16_SLV_LEN-1 downto 0);
  begin

        data_slv := data((pos+uint32_t_16_SLV_LEN)-1 downto pos);
        rv.data := slv_to_uint32_t_16(data_slv);
        pos := pos + uint32_t_16_SLV_LEN;

      return rv;
  end function;

  function uint8_t_array_144_t_to_slv(data : uint8_t_array_144_t) return std_logic_vector is
    variable rv : std_logic_vector(uint8_t_array_144_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+uint8_t_144_SLV_LEN)-1 downto pos) := uint8_t_144_to_slv(data.data);
        pos := pos + uint8_t_144_SLV_LEN;

      return rv;
  end function;

  function slv_to_uint8_t_array_144_t(data : std_logic_vector) return uint8_t_array_144_t is
    variable rv : uint8_t_array_144_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(uint8_t_144_SLV_LEN-1 downto 0);
  begin

        data_slv := data((pos+uint8_t_144_SLV_LEN)-1 downto pos);
        rv.data := slv_to_uint8_t_144(data_slv);
        pos := pos + uint8_t_144_SLV_LEN;

      return rv;
  end function;

  function char_array_128_t_to_slv(data : char_array_128_t) return std_logic_vector is
    variable rv : std_logic_vector(char_array_128_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+char_128_SLV_LEN)-1 downto pos) := char_128_to_slv(data.data);
        pos := pos + char_128_SLV_LEN;

      return rv;
  end function;

  function slv_to_char_array_128_t(data : std_logic_vector) return char_array_128_t is
    variable rv : char_array_128_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(char_128_SLV_LEN-1 downto 0);
  begin

        data_slv := data((pos+char_128_SLV_LEN)-1 downto pos);
        rv.data := slv_to_char_128(data_slv);
        pos := pos + char_128_SLV_LEN;

      return rv;
  end function;

      function axis128_t_stream_t_4_to_slv(data : axis128_t_stream_t_4) return std_logic_vector is
        variable rv : std_logic_vector(axis128_t_stream_t_4_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos) := axis128_t_stream_t_to_slv(data(0));
            pos := pos + axis128_t_stream_t_SLV_LEN;
    
            rv((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos) := axis128_t_stream_t_to_slv(data(1));
            pos := pos + axis128_t_stream_t_SLV_LEN;
    
            rv((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos) := axis128_t_stream_t_to_slv(data(2));
            pos := pos + axis128_t_stream_t_SLV_LEN;
    
            rv((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos) := axis128_t_stream_t_to_slv(data(3));
            pos := pos + axis128_t_stream_t_SLV_LEN;
    
          return rv;
      end function;
    
      function slv_to_axis128_t_stream_t_4(data : std_logic_vector) return axis128_t_stream_t_4 is
        variable rv : axis128_t_stream_t_4;
        variable elem_slv : std_logic_vector(axis128_t_stream_t_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos);
            rv(0) := slv_to_axis128_t_stream_t(elem_slv);
            pos := pos + axis128_t_stream_t_SLV_LEN;
    
            elem_slv := data((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos);
            rv(1) := slv_to_axis128_t_stream_t(elem_slv);
            pos := pos + axis128_t_stream_t_SLV_LEN;
    
            elem_slv := data((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos);
            rv(2) := slv_to_axis128_t_stream_t(elem_slv);
            pos := pos + axis128_t_stream_t_SLV_LEN;
    
            elem_slv := data((pos+axis128_t_stream_t_SLV_LEN)-1 downto pos);
            rv(3) := slv_to_axis128_t_stream_t(elem_slv);
            pos := pos + axis128_t_stream_t_SLV_LEN;
    
          return rv;
      end function;
    
      function axis128_t_1_to_slv(data : axis128_t_1) return std_logic_vector is
        variable rv : std_logic_vector(axis128_t_1_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            rv((pos+axis128_t_SLV_LEN)-1 downto pos) := axis128_t_to_slv(data(0));
            pos := pos + axis128_t_SLV_LEN;
    
          return rv;
      end function;
    
      function slv_to_axis128_t_1(data : std_logic_vector) return axis128_t_1 is
        variable rv : axis128_t_1;
        variable elem_slv : std_logic_vector(axis128_t_SLV_LEN-1 downto 0);
        variable pos : integer := 0;
      begin
    
            elem_slv := data((pos+axis128_t_SLV_LEN)-1 downto pos);
            rv(0) := slv_to_axis128_t(elem_slv);
            pos := pos + axis128_t_SLV_LEN;
    
          return rv;
      end function;
    
  function axis512_to_axis128_array_t_to_slv(data : axis512_to_axis128_array_t) return std_logic_vector is
    variable rv : std_logic_vector(axis512_to_axis128_array_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis128_t_stream_t_4_SLV_LEN)-1 downto pos) := axis128_t_stream_t_4_to_slv(data.axis_chunks);
        pos := pos + axis128_t_stream_t_4_SLV_LEN;

      return rv;
  end function;

  function slv_to_axis512_to_axis128_array_t(data : std_logic_vector) return axis512_to_axis128_array_t is
    variable rv : axis512_to_axis128_array_t;
    variable pos : integer := 0;
    variable axis_chunks_slv : std_logic_vector(axis128_t_stream_t_4_SLV_LEN-1 downto 0);
  begin

        axis_chunks_slv := data((pos+axis128_t_stream_t_4_SLV_LEN)-1 downto pos);
        rv.axis_chunks := slv_to_axis128_t_stream_t_4(axis_chunks_slv);
        pos := pos + axis128_t_stream_t_4_SLV_LEN;

      return rv;
  end function;

  function verify_fifo_FIFO_read_t_to_slv(data : verify_fifo_FIFO_read_t) return std_logic_vector is
    variable rv : std_logic_vector(verify_fifo_FIFO_read_t_SLV_LEN-1 downto 0);
    variable pos : integer := 0;
  begin

        rv((pos+axis128_t_1_SLV_LEN)-1 downto pos) := axis128_t_1_to_slv(data.data);
        pos := pos + axis128_t_1_SLV_LEN;

        rv((pos+1)-1 downto pos) := std_logic_vector(data.valid);
        pos := pos + 1;

      return rv;
  end function;

  function slv_to_verify_fifo_FIFO_read_t(data : std_logic_vector) return verify_fifo_FIFO_read_t is
    variable rv : verify_fifo_FIFO_read_t;
    variable pos : integer := 0;
    variable data_slv : std_logic_vector(axis128_t_1_SLV_LEN-1 downto 0);
    variable valid_slv : std_logic_vector(1-1 downto 0);
  begin

        data_slv := data((pos+axis128_t_1_SLV_LEN)-1 downto pos);
        rv.data := slv_to_axis128_t_1(data_slv);
        pos := pos + axis128_t_1_SLV_LEN;

        valid_slv := data((pos+1)-1 downto pos);
        rv.valid := unsigned(valid_slv);
        pos := pos + 1;

      return rv;
  end function;
end package body c_structs_pkg;
