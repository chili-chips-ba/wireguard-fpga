mem['h0000] = 32'h00001517;
mem['h0001] = 32'h25850513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'h00860613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFE850513;
mem['h000E] = 32'h10001597;
mem['h000F] = 32'h3F458593;
mem['h0010] = 32'h00B55863;
mem['h0011] = 32'h00052023;
mem['h0012] = 32'h00450513;
mem['h0013] = 32'hFEB54CE3;
mem['h0014] = 32'h10008117;
mem['h0015] = 32'hFB010113;
mem['h0016] = 32'h10000197;
mem['h0017] = 32'h7C018193;
mem['h0018] = 32'h00A54533;
mem['h0019] = 32'h00B5C5B3;
mem['h001A] = 32'h00C64633;
mem['h001B] = 32'h518000EF;
mem['h001C] = 32'h0000006F;
mem['h001D] = 32'h00452783;
mem['h001E] = 32'h0087A783;
mem['h001F] = 32'h0007A783;
mem['h0020] = 32'h0007A783;
mem['h0021] = 32'hFE07C8E3;
mem['h0022] = 32'h00452783;
mem['h0023] = 32'h0087A783;
mem['h0024] = 32'h0007A783;
mem['h0025] = 32'h00B78023;
mem['h0026] = 32'h00008067;
mem['h0027] = 32'h0A058A63;
mem['h0028] = 32'hFE010113;
mem['h0029] = 32'h00912A23;
mem['h002A] = 32'h00058493;
mem['h002B] = 32'h01212823;
mem['h002C] = 32'h00A00593;
mem['h002D] = 32'h00050913;
mem['h002E] = 32'h00048513;
mem['h002F] = 32'h00812C23;
mem['h0030] = 32'h00112E23;
mem['h0031] = 32'h01312623;
mem['h0032] = 32'h01412423;
mem['h0033] = 32'h729000EF;
mem['h0034] = 32'h01051513;
mem['h0035] = 32'h01055513;
mem['h0036] = 32'h00100413;
mem['h0037] = 32'h06857E63;
mem['h0038] = 32'h00900A13;
mem['h0039] = 32'h00040593;
mem['h003A] = 32'h00048513;
mem['h003B] = 32'h709000EF;
mem['h003C] = 32'h03050593;
mem['h003D] = 32'h0FF5F593;
mem['h003E] = 32'h00090513;
mem['h003F] = 32'hF79FF0EF;
mem['h0040] = 32'h00040593;
mem['h0041] = 32'h00048513;
mem['h0042] = 32'h735000EF;
mem['h0043] = 32'h01051493;
mem['h0044] = 32'h00A00593;
mem['h0045] = 32'h00040513;
mem['h0046] = 32'h6DD000EF;
mem['h0047] = 32'h00040993;
mem['h0048] = 32'h01051413;
mem['h0049] = 32'h0104D493;
mem['h004A] = 32'h01045413;
mem['h004B] = 32'hFB3A6CE3;
mem['h004C] = 32'h01C12083;
mem['h004D] = 32'h01812403;
mem['h004E] = 32'h01412483;
mem['h004F] = 32'h01012903;
mem['h0050] = 32'h00C12983;
mem['h0051] = 32'h00812A03;
mem['h0052] = 32'h02010113;
mem['h0053] = 32'h00008067;
mem['h0054] = 32'h03000593;
mem['h0055] = 32'hF21FF06F;
mem['h0056] = 32'h00241793;
mem['h0057] = 32'h00F40433;
mem['h0058] = 32'h00141413;
mem['h0059] = 32'h01041413;
mem['h005A] = 32'h01045413;
mem['h005B] = 32'hF71FF06F;
mem['h005C] = 32'hFF010113;
mem['h005D] = 32'h00812423;
mem['h005E] = 32'h00912223;
mem['h005F] = 32'h00112623;
mem['h0060] = 32'h00050493;
mem['h0061] = 32'h00058413;
mem['h0062] = 32'h00044583;
mem['h0063] = 32'h00059C63;
mem['h0064] = 32'h00C12083;
mem['h0065] = 32'h00812403;
mem['h0066] = 32'h00412483;
mem['h0067] = 32'h01010113;
mem['h0068] = 32'h00008067;
mem['h0069] = 32'h00048513;
mem['h006A] = 32'h00140413;
mem['h006B] = 32'hEC9FF0EF;
mem['h006C] = 32'hFD9FF06F;
mem['h006D] = 32'hFF010113;
mem['h006E] = 32'h00112623;
mem['h006F] = 32'h00812423;
mem['h0070] = 32'h00912223;
mem['h0071] = 32'h00058493;
mem['h0072] = 32'h0005C583;
mem['h0073] = 32'h00050413;
mem['h0074] = 32'hECDFF0EF;
mem['h0075] = 32'h00040513;
mem['h0076] = 32'h02E00593;
mem['h0077] = 32'hE99FF0EF;
mem['h0078] = 32'h0014C583;
mem['h0079] = 32'h00040513;
mem['h007A] = 32'hEB5FF0EF;
mem['h007B] = 32'h00040513;
mem['h007C] = 32'h02E00593;
mem['h007D] = 32'hE81FF0EF;
mem['h007E] = 32'h0024C583;
mem['h007F] = 32'h00040513;
mem['h0080] = 32'hE9DFF0EF;
mem['h0081] = 32'h00040513;
mem['h0082] = 32'h02E00593;
mem['h0083] = 32'hE69FF0EF;
mem['h0084] = 32'h00040513;
mem['h0085] = 32'h00812403;
mem['h0086] = 32'h0034C583;
mem['h0087] = 32'h00C12083;
mem['h0088] = 32'h00412483;
mem['h0089] = 32'h01010113;
mem['h008A] = 32'hE75FF06F;
mem['h008B] = 32'h00100613;
mem['h008C] = 32'h00010837;
mem['h008D] = 32'h00050693;
mem['h008E] = 32'h00000793;
mem['h008F] = 32'h40A60633;
mem['h0090] = 32'hFFF80893;
mem['h0091] = 32'h00D60733;
mem['h0092] = 32'h04B76063;
mem['h0093] = 32'hFFE5F713;
mem['h0094] = 32'h02B77463;
mem['h0095] = 32'h00E50533;
mem['h0096] = 32'h00054703;
mem['h0097] = 32'h00871713;
mem['h0098] = 32'h00E787B3;
mem['h0099] = 32'h00010737;
mem['h009A] = 32'h00E7E863;
mem['h009B] = 32'h01079793;
mem['h009C] = 32'h0107D793;
mem['h009D] = 32'h00178793;
mem['h009E] = 32'hFFF7C513;
mem['h009F] = 32'h01051513;
mem['h00A0] = 32'h01055513;
mem['h00A1] = 32'h00008067;
mem['h00A2] = 32'h0006C703;
mem['h00A3] = 32'h0016C303;
mem['h00A4] = 32'h00871713;
mem['h00A5] = 32'h00676733;
mem['h00A6] = 32'h01071713;
mem['h00A7] = 32'h01075713;
mem['h00A8] = 32'h00E787B3;
mem['h00A9] = 32'h0107E663;
mem['h00AA] = 32'h0117F7B3;
mem['h00AB] = 32'h00178793;
mem['h00AC] = 32'h00268693;
mem['h00AD] = 32'hF91FF06F;
mem['h00AE] = 32'h100016B7;
mem['h00AF] = 32'h4286A703;
mem['h00B0] = 32'h100017B7;
mem['h00B1] = 32'hC2878793;
mem['h00B2] = 32'h00F707B3;
mem['h00B3] = 32'h00A70733;
mem['h00B4] = 32'h42E6A423;
mem['h00B5] = 32'h000016B7;
mem['h00B6] = 32'h80068693;
mem['h00B7] = 32'h00E6D463;
mem['h00B8] = 32'h00100073;
mem['h00B9] = 32'h00078513;
mem['h00BA] = 32'h00008067;
mem['h00BB] = 32'hFF010113;
mem['h00BC] = 32'h00812423;
mem['h00BD] = 32'h00001437;
mem['h00BE] = 32'h0A040413;
mem['h00BF] = 32'h0045D793;
mem['h00C0] = 32'h00F407B3;
mem['h00C1] = 32'h00912223;
mem['h00C2] = 32'h00058493;
mem['h00C3] = 32'h0007C583;
mem['h00C4] = 32'h00F4F493;
mem['h00C5] = 32'h01212023;
mem['h00C6] = 32'h00112623;
mem['h00C7] = 32'h00050913;
mem['h00C8] = 32'h00940433;
mem['h00C9] = 32'hD51FF0EF;
mem['h00CA] = 32'h00044583;
mem['h00CB] = 32'h00812403;
mem['h00CC] = 32'h00C12083;
mem['h00CD] = 32'h00412483;
mem['h00CE] = 32'h00090513;
mem['h00CF] = 32'h00012903;
mem['h00D0] = 32'h01010113;
mem['h00D1] = 32'hD31FF06F;
mem['h00D2] = 32'h00000793;
mem['h00D3] = 32'h00C79463;
mem['h00D4] = 32'h00008067;
mem['h00D5] = 32'h00F58733;
mem['h00D6] = 32'h00074683;
mem['h00D7] = 32'h00F50733;
mem['h00D8] = 32'h00178793;
mem['h00D9] = 32'h00D70023;
mem['h00DA] = 32'hFE5FF06F;
mem['h00DB] = 32'h00052783;
mem['h00DC] = 32'h0007A783;
mem['h00DD] = 32'h0187A783;
mem['h00DE] = 32'h0007A783;
mem['h00DF] = 32'h0007A783;
mem['h00E0] = 32'h0017F793;
mem['h00E1] = 32'h1E078E63;
mem['h00E2] = 32'h00052783;
mem['h00E3] = 32'h0005C703;
mem['h00E4] = 32'hFFFF8637;
mem['h00E5] = 32'h0007A783;
mem['h00E6] = 32'h00777713;
mem['h00E7] = 32'hFFFF08B7;
mem['h00E8] = 32'h0107A783;
mem['h00E9] = 32'hFFF60613;
mem['h00EA] = 32'h0007A683;
mem['h00EB] = 32'h0006A783;
mem['h00EC] = 32'hFF87F793;
mem['h00ED] = 32'h00E7E7B3;
mem['h00EE] = 32'h00F6A023;
mem['h00EF] = 32'h00052783;
mem['h00F0] = 32'h0015C703;
mem['h00F1] = 32'h0007A783;
mem['h00F2] = 32'h00777713;
mem['h00F3] = 32'h00371713;
mem['h00F4] = 32'h0107A783;
mem['h00F5] = 32'h0007A683;
mem['h00F6] = 32'h0006A783;
mem['h00F7] = 32'hFC77F793;
mem['h00F8] = 32'h00E7E7B3;
mem['h00F9] = 32'h00F6A023;
mem['h00FA] = 32'h00052783;
mem['h00FB] = 32'h0025C703;
mem['h00FC] = 32'h0007A783;
mem['h00FD] = 32'h00177713;
mem['h00FE] = 32'h00671713;
mem['h00FF] = 32'h0107A783;
mem['h0100] = 32'h0007A683;
mem['h0101] = 32'h0006A783;
mem['h0102] = 32'hFBF7F793;
mem['h0103] = 32'h00E7E7B3;
mem['h0104] = 32'h00F6A023;
mem['h0105] = 32'h00052783;
mem['h0106] = 32'h0035C703;
mem['h0107] = 32'h0007A783;
mem['h0108] = 32'h00177713;
mem['h0109] = 32'h00771713;
mem['h010A] = 32'h0107A783;
mem['h010B] = 32'h0007A683;
mem['h010C] = 32'h0006A783;
mem['h010D] = 32'hF7F7F793;
mem['h010E] = 32'h00E7E7B3;
mem['h010F] = 32'h00F6A023;
mem['h0110] = 32'h00858713;
mem['h0111] = 32'h00000793;
mem['h0112] = 32'h00052683;
mem['h0113] = 32'h00072803;
mem['h0114] = 32'h01078793;
mem['h0115] = 32'h0006A683;
mem['h0116] = 32'h01070713;
mem['h0117] = 32'h0006A683;
mem['h0118] = 32'h0006A683;
mem['h0119] = 32'h0106A023;
mem['h011A] = 32'h00052683;
mem['h011B] = 32'hFF472803;
mem['h011C] = 32'h0006A683;
mem['h011D] = 32'h0046A683;
mem['h011E] = 32'h0006A683;
mem['h011F] = 32'h0106A023;
mem['h0120] = 32'h00052683;
mem['h0121] = 32'hFF872803;
mem['h0122] = 32'h0006A683;
mem['h0123] = 32'h0086A683;
mem['h0124] = 32'h0006A683;
mem['h0125] = 32'h0106A023;
mem['h0126] = 32'h00052683;
mem['h0127] = 32'hFFC72803;
mem['h0128] = 32'h0006A683;
mem['h0129] = 32'h00C6A683;
mem['h012A] = 32'h0006A683;
mem['h012B] = 32'h0106A023;
mem['h012C] = 32'h0045A683;
mem['h012D] = 32'h04D7FE63;
mem['h012E] = 32'h00052683;
mem['h012F] = 32'h0006A683;
mem['h0130] = 32'h0106A683;
mem['h0131] = 32'h0006A803;
mem['h0132] = 32'h00082683;
mem['h0133] = 32'h0116E6B3;
mem['h0134] = 32'h00D82023;
mem['h0135] = 32'h00052683;
mem['h0136] = 32'h0006A683;
mem['h0137] = 32'h0106A683;
mem['h0138] = 32'h0006A803;
mem['h0139] = 32'h00082683;
mem['h013A] = 32'h00C6F6B3;
mem['h013B] = 32'h00D82023;
mem['h013C] = 32'h00052683;
mem['h013D] = 32'h0006A683;
mem['h013E] = 32'h0146A683;
mem['h013F] = 32'h0006A803;
mem['h0140] = 32'h00082683;
mem['h0141] = 32'h0016E693;
mem['h0142] = 32'h00D82023;
mem['h0143] = 32'hF3DFF06F;
mem['h0144] = 32'h00052703;
mem['h0145] = 32'h40D787B3;
mem['h0146] = 32'h000106B7;
mem['h0147] = 32'h00072703;
mem['h0148] = 32'hFFF68693;
mem['h0149] = 32'h40F6D7B3;
mem['h014A] = 32'h01072703;
mem['h014B] = 32'h01079793;
mem['h014C] = 32'h00072603;
mem['h014D] = 32'h00062703;
mem['h014E] = 32'h00D77733;
mem['h014F] = 32'h00F767B3;
mem['h0150] = 32'h00F62023;
mem['h0151] = 32'h00052783;
mem['h0152] = 32'h000086B7;
mem['h0153] = 32'h0007A783;
mem['h0154] = 32'h0107A783;
mem['h0155] = 32'h0007A703;
mem['h0156] = 32'h00072783;
mem['h0157] = 32'h00D7E7B3;
mem['h0158] = 32'h00F72023;
mem['h0159] = 32'h00052783;
mem['h015A] = 32'h0007A783;
mem['h015B] = 32'h0147A783;
mem['h015C] = 32'h0007A703;
mem['h015D] = 32'h00072783;
mem['h015E] = 32'h0017E793;
mem['h015F] = 32'h00F72023;
mem['h0160] = 32'h00008067;
mem['h0161] = 32'hF9010113;
mem['h0162] = 32'h02400513;
mem['h0163] = 32'h06112623;
mem['h0164] = 32'h06812423;
mem['h0165] = 32'h06912223;
mem['h0166] = 32'h07212023;
mem['h0167] = 32'h05312E23;
mem['h0168] = 32'h05412C23;
mem['h0169] = 32'h05512A23;
mem['h016A] = 32'h05612823;
mem['h016B] = 32'h05712623;
mem['h016C] = 32'h05812423;
mem['h016D] = 32'h05912223;
mem['h016E] = 32'h05A12023;
mem['h016F] = 32'h03B12E23;
mem['h0170] = 32'hCF9FF0EF;
mem['h0171] = 32'h00050413;
mem['h0172] = 32'h00800513;
mem['h0173] = 32'hCEDFF0EF;
mem['h0174] = 32'h00050913;
mem['h0175] = 32'h01C00513;
mem['h0176] = 32'hCE1FF0EF;
mem['h0177] = 32'h00050493;
mem['h0178] = 32'h00400513;
mem['h0179] = 32'hCD5FF0EF;
mem['h017A] = 32'h200007B7;
mem['h017B] = 32'h00F52023;
mem['h017C] = 32'h00A4A023;
mem['h017D] = 32'h00400513;
mem['h017E] = 32'hCC1FF0EF;
mem['h017F] = 32'h200007B7;
mem['h0180] = 32'h00478793;
mem['h0181] = 32'h00F52023;
mem['h0182] = 32'h00A4A223;
mem['h0183] = 32'h00400513;
mem['h0184] = 32'hCA9FF0EF;
mem['h0185] = 32'h200007B7;
mem['h0186] = 32'h00878793;
mem['h0187] = 32'h00F52023;
mem['h0188] = 32'h00A4A423;
mem['h0189] = 32'h00400513;
mem['h018A] = 32'hC91FF0EF;
mem['h018B] = 32'h200007B7;
mem['h018C] = 32'h00C78793;
mem['h018D] = 32'h00F52023;
mem['h018E] = 32'h00A4A623;
mem['h018F] = 32'h00400513;
mem['h0190] = 32'hC79FF0EF;
mem['h0191] = 32'h200007B7;
mem['h0192] = 32'h01078793;
mem['h0193] = 32'h00F52023;
mem['h0194] = 32'h00A4A823;
mem['h0195] = 32'h00400513;
mem['h0196] = 32'hC61FF0EF;
mem['h0197] = 32'h200007B7;
mem['h0198] = 32'h01478793;
mem['h0199] = 32'h00F52023;
mem['h019A] = 32'h00A4AA23;
mem['h019B] = 32'h00400513;
mem['h019C] = 32'hC49FF0EF;
mem['h019D] = 32'h200007B7;
mem['h019E] = 32'h01878793;
mem['h019F] = 32'h00F52023;
mem['h01A0] = 32'h00A4AC23;
mem['h01A1] = 32'h00992023;
mem['h01A2] = 32'h01C00513;
mem['h01A3] = 32'hC2DFF0EF;
mem['h01A4] = 32'h00050493;
mem['h01A5] = 32'h00400513;
mem['h01A6] = 32'hC21FF0EF;
mem['h01A7] = 32'h200007B7;
mem['h01A8] = 32'h01C78793;
mem['h01A9] = 32'h00F52023;
mem['h01AA] = 32'h00A4A023;
mem['h01AB] = 32'h00400513;
mem['h01AC] = 32'hC09FF0EF;
mem['h01AD] = 32'h200007B7;
mem['h01AE] = 32'h02078793;
mem['h01AF] = 32'h00F52023;
mem['h01B0] = 32'h00A4A223;
mem['h01B1] = 32'h00400513;
mem['h01B2] = 32'hBF1FF0EF;
mem['h01B3] = 32'h200007B7;
mem['h01B4] = 32'h02478793;
mem['h01B5] = 32'h00F52023;
mem['h01B6] = 32'h00A4A423;
mem['h01B7] = 32'h00400513;
mem['h01B8] = 32'hBD9FF0EF;
mem['h01B9] = 32'h200007B7;
mem['h01BA] = 32'h02878793;
mem['h01BB] = 32'h00F52023;
mem['h01BC] = 32'h00A4A623;
mem['h01BD] = 32'h00400513;
mem['h01BE] = 32'hBC1FF0EF;
mem['h01BF] = 32'h200007B7;
mem['h01C0] = 32'h02C78793;
mem['h01C1] = 32'h00F52023;
mem['h01C2] = 32'h00A4A823;
mem['h01C3] = 32'h00400513;
mem['h01C4] = 32'hBA9FF0EF;
mem['h01C5] = 32'h200007B7;
mem['h01C6] = 32'h03078793;
mem['h01C7] = 32'h00F52023;
mem['h01C8] = 32'h00A4AA23;
mem['h01C9] = 32'h00400513;
mem['h01CA] = 32'hB91FF0EF;
mem['h01CB] = 32'h200007B7;
mem['h01CC] = 32'h03478793;
mem['h01CD] = 32'h00F52023;
mem['h01CE] = 32'h00A4AC23;
mem['h01CF] = 32'h00992223;
mem['h01D0] = 32'h01242023;
mem['h01D1] = 32'h01000513;
mem['h01D2] = 32'hB71FF0EF;
mem['h01D3] = 32'h00050493;
mem['h01D4] = 32'h00400513;
mem['h01D5] = 32'hB65FF0EF;
mem['h01D6] = 32'h200007B7;
mem['h01D7] = 32'h03878793;
mem['h01D8] = 32'h00F52023;
mem['h01D9] = 32'h00A4A023;
mem['h01DA] = 32'h00400513;
mem['h01DB] = 32'hB4DFF0EF;
mem['h01DC] = 32'h200007B7;
mem['h01DD] = 32'h03C78793;
mem['h01DE] = 32'h00F52023;
mem['h01DF] = 32'h00A4A223;
mem['h01E0] = 32'h00400513;
mem['h01E1] = 32'hB35FF0EF;
mem['h01E2] = 32'h200007B7;
mem['h01E3] = 32'h04078793;
mem['h01E4] = 32'h00F52023;
mem['h01E5] = 32'h00A4A423;
mem['h01E6] = 32'h00400513;
mem['h01E7] = 32'hB1DFF0EF;
mem['h01E8] = 32'h200007B7;
mem['h01E9] = 32'h04478793;
mem['h01EA] = 32'h00F52023;
mem['h01EB] = 32'h00A4A623;
mem['h01EC] = 32'h00942223;
mem['h01ED] = 32'h00400513;
mem['h01EE] = 32'hB01FF0EF;
mem['h01EF] = 32'h200007B7;
mem['h01F0] = 32'h04878793;
mem['h01F1] = 32'h00F52023;
mem['h01F2] = 32'h200004B7;
mem['h01F3] = 32'hE0000A37;
mem['h01F4] = 32'h200009B7;
mem['h01F5] = 32'h00A42423;
mem['h01F6] = 32'h04C48493;
mem['h01F7] = 32'hFC0A0A13;
mem['h01F8] = 32'h05C98993;
mem['h01F9] = 32'h00400513;
mem['h01FA] = 32'hAD1FF0EF;
mem['h01FB] = 32'h00050913;
mem['h01FC] = 32'h00400513;
mem['h01FD] = 32'hAC5FF0EF;
mem['h01FE] = 32'h00952023;
mem['h01FF] = 32'h014487B3;
mem['h0200] = 32'h00A92023;
mem['h0201] = 32'h00F407B3;
mem['h0202] = 32'h0127A023;
mem['h0203] = 32'h00448493;
mem['h0204] = 32'hFD349AE3;
mem['h0205] = 32'h00400513;
mem['h0206] = 32'hAA1FF0EF;
mem['h0207] = 32'h00050913;
mem['h0208] = 32'h00400513;
mem['h0209] = 32'hA95FF0EF;
mem['h020A] = 32'h00952023;
mem['h020B] = 32'h00A92023;
mem['h020C] = 32'h01242E23;
mem['h020D] = 32'h00400513;
mem['h020E] = 32'hA81FF0EF;
mem['h020F] = 32'h200007B7;
mem['h0210] = 32'h06078793;
mem['h0211] = 32'h00F52023;
mem['h0212] = 32'h000014B7;
mem['h0213] = 32'h0B448593;
mem['h0214] = 32'h02A42023;
mem['h0215] = 32'h00040513;
mem['h0216] = 32'h919FF0EF;
mem['h0217] = 32'h000015B7;
mem['h0218] = 32'h0E458593;
mem['h0219] = 32'h00040513;
mem['h021A] = 32'h909FF0EF;
mem['h021B] = 32'h0B448593;
mem['h021C] = 32'h00040513;
mem['h021D] = 32'h8FDFF0EF;
mem['h021E] = 32'h000015B7;
mem['h021F] = 32'h11458593;
mem['h0220] = 32'h00040513;
mem['h0221] = 32'h8EDFF0EF;
mem['h0222] = 32'h000015B7;
mem['h0223] = 32'h12C58593;
mem['h0224] = 32'h00040513;
mem['h0225] = 32'h8DDFF0EF;
mem['h0226] = 32'h10000937;
mem['h0227] = 32'h00090593;
mem['h0228] = 32'h00040513;
mem['h0229] = 32'h911FF0EF;
mem['h022A] = 32'h000015B7;
mem['h022B] = 32'h14458593;
mem['h022C] = 32'h00040513;
mem['h022D] = 32'h00090493;
mem['h022E] = 32'h8B9FF0EF;
mem['h022F] = 32'h00448593;
mem['h0230] = 32'h00040513;
mem['h0231] = 32'h8F1FF0EF;
mem['h0232] = 32'h000015B7;
mem['h0233] = 32'h16058593;
mem['h0234] = 32'h00040513;
mem['h0235] = 32'h89DFF0EF;
mem['h0236] = 32'h0084C583;
mem['h0237] = 32'h00040513;
mem['h0238] = 32'h100009B7;
mem['h0239] = 32'hA09FF0EF;
mem['h023A] = 32'h03A00593;
mem['h023B] = 32'h00040513;
mem['h023C] = 32'hF84FF0EF;
mem['h023D] = 32'h0094C583;
mem['h023E] = 32'h00040513;
mem['h023F] = 32'h01898A93;
mem['h0240] = 32'h9EDFF0EF;
mem['h0241] = 32'h03A00593;
mem['h0242] = 32'h00040513;
mem['h0243] = 32'hF68FF0EF;
mem['h0244] = 32'h00A4C583;
mem['h0245] = 32'h00040513;
mem['h0246] = 32'h00090A13;
mem['h0247] = 32'h9D1FF0EF;
mem['h0248] = 32'h03A00593;
mem['h0249] = 32'h00040513;
mem['h024A] = 32'hF4CFF0EF;
mem['h024B] = 32'h00B4C583;
mem['h024C] = 32'h00040513;
mem['h024D] = 32'h9B9FF0EF;
mem['h024E] = 32'h03A00593;
mem['h024F] = 32'h00040513;
mem['h0250] = 32'hF34FF0EF;
mem['h0251] = 32'h00C4C583;
mem['h0252] = 32'h00040513;
mem['h0253] = 32'h9A1FF0EF;
mem['h0254] = 32'h03A00593;
mem['h0255] = 32'h00040513;
mem['h0256] = 32'hF1CFF0EF;
mem['h0257] = 32'h00D4C583;
mem['h0258] = 32'h00040513;
mem['h0259] = 32'h989FF0EF;
mem['h025A] = 32'h000015B7;
mem['h025B] = 32'h17C58593;
mem['h025C] = 32'h00040513;
mem['h025D] = 32'hFFCFF0EF;
mem['h025E] = 32'h00E48593;
mem['h025F] = 32'h00040513;
mem['h0260] = 32'h835FF0EF;
mem['h0261] = 32'h000015B7;
mem['h0262] = 32'h19858593;
mem['h0263] = 32'h00040513;
mem['h0264] = 32'hFE0FF0EF;
mem['h0265] = 32'h0124C583;
mem['h0266] = 32'h00040513;
mem['h0267] = 32'h000014B7;
mem['h0268] = 32'hEFCFF0EF;
mem['h0269] = 32'h1B448593;
mem['h026A] = 32'h00040513;
mem['h026B] = 32'hFC4FF0EF;
mem['h026C] = 32'h000015B7;
mem['h026D] = 32'h1B858593;
mem['h026E] = 32'h00040513;
mem['h026F] = 32'hFB4FF0EF;
mem['h0270] = 32'h608A8793;
mem['h0271] = 32'h00F12423;
mem['h0272] = 32'h00F12623;
mem['h0273] = 32'h00A00B13;
mem['h0274] = 32'h00D00B93;
mem['h0275] = 32'h000A8023;
mem['h0276] = 32'h000A9123;
mem['h0277] = 32'h00042703;
mem['h0278] = 32'h00472703;
mem['h0279] = 32'h01872703;
mem['h027A] = 32'h00072703;
mem['h027B] = 32'h00072703;
mem['h027C] = 32'h00177713;
mem['h027D] = 32'h10070463;
mem['h027E] = 32'h00042703;
mem['h027F] = 32'h000A8C93;
mem['h0280] = 32'h01898693;
mem['h0281] = 32'h00472703;
mem['h0282] = 32'h5F000513;
mem['h0283] = 32'h01072703;
mem['h0284] = 32'h00072703;
mem['h0285] = 32'h00072703;
mem['h0286] = 32'h00375713;
mem['h0287] = 32'h00777713;
mem['h0288] = 32'h00EA80A3;
mem['h0289] = 32'h00000713;
mem['h028A] = 32'h06E56263;
mem['h028B] = 32'h00042603;
mem['h028C] = 32'h00462603;
mem['h028D] = 32'h00062603;
mem['h028E] = 32'h00062603;
mem['h028F] = 32'h00062603;
mem['h0290] = 32'h00C6A423;
mem['h0291] = 32'h00042603;
mem['h0292] = 32'h00462603;
mem['h0293] = 32'h00462603;
mem['h0294] = 32'h00062603;
mem['h0295] = 32'h00062603;
mem['h0296] = 32'h00C6A623;
mem['h0297] = 32'h00042603;
mem['h0298] = 32'h00462603;
mem['h0299] = 32'h00862603;
mem['h029A] = 32'h00062603;
mem['h029B] = 32'h00062603;
mem['h029C] = 32'h00C6A823;
mem['h029D] = 32'h00042603;
mem['h029E] = 32'h00462603;
mem['h029F] = 32'h00C62603;
mem['h02A0] = 32'h00062603;
mem['h02A1] = 32'h00062603;
mem['h02A2] = 32'h00C6AA23;
mem['h02A3] = 32'h00042603;
mem['h02A4] = 32'h01068693;
mem['h02A5] = 32'h00462603;
mem['h02A6] = 32'h01062603;
mem['h02A7] = 32'h00062603;
mem['h02A8] = 32'h00062603;
mem['h02A9] = 32'h01061593;
mem['h02AA] = 32'h0605DC63;
mem['h02AB] = 32'h00042683;
mem['h02AC] = 32'h0046A683;
mem['h02AD] = 32'h0106A683;
mem['h02AE] = 32'h0006A683;
mem['h02AF] = 32'h0026D683;
mem['h02B0] = 32'h0016F613;
mem['h02B1] = 32'h04061863;
mem['h02B2] = 32'h60000693;
mem['h02B3] = 32'h00E6F463;
mem['h02B4] = 32'h60000713;
mem['h02B5] = 32'h00EAA223;
mem['h02B6] = 32'h00042703;
mem['h02B7] = 32'h00472703;
mem['h02B8] = 32'h01472703;
mem['h02B9] = 32'h00072683;
mem['h02BA] = 32'h0006A703;
mem['h02BB] = 32'h00176713;
mem['h02BC] = 32'h00E6A023;
mem['h02BD] = 32'h004AA703;
mem['h02BE] = 32'h04071663;
mem['h02BF] = 32'h00842703;
mem['h02C0] = 32'h00072683;
mem['h02C1] = 32'h0006A703;
mem['h02C2] = 32'hDFF77713;
mem['h02C3] = 32'h00E6A023;
mem['h02C4] = 32'h3500006F;
mem['h02C5] = 32'h00170713;
mem['h02C6] = 32'h0016D693;
mem['h02C7] = 32'hFA5FF06F;
mem['h02C8] = 32'h00042603;
mem['h02C9] = 32'h01070713;
mem['h02CA] = 32'h00462603;
mem['h02CB] = 32'h01462603;
mem['h02CC] = 32'h00062583;
mem['h02CD] = 32'h0005A603;
mem['h02CE] = 32'h00166613;
mem['h02CF] = 32'h00C5A023;
mem['h02D0] = 32'hEE9FF06F;
mem['h02D1] = 32'h00842703;
mem['h02D2] = 32'h00072683;
mem['h02D3] = 32'h0006A703;
mem['h02D4] = 32'h20076713;
mem['h02D5] = 32'h00E6A023;
mem['h02D6] = 32'h014ACD03;
mem['h02D7] = 32'h00800713;
mem['h02D8] = 32'h2CED1E63;
mem['h02D9] = 32'h015AC703;
mem['h02DA] = 32'h00600693;
mem['h02DB] = 32'h18D70263;
mem['h02DC] = 32'h2C071663;
mem['h02DD] = 32'h016AC703;
mem['h02DE] = 32'h04000693;
mem['h02DF] = 32'h0F077713;
mem['h02E0] = 32'h2AD71E63;
mem['h02E1] = 32'h01FAC683;
mem['h02E2] = 32'h00100713;
mem['h02E3] = 32'h2AE69863;
mem['h02E4] = 32'h000015B7;
mem['h02E5] = 32'h1E858593;
mem['h02E6] = 32'h00040513;
mem['h02E7] = 32'hDD4FF0EF;
mem['h02E8] = 32'h004AD583;
mem['h02E9] = 32'h00040513;
mem['h02EA] = 32'hCF4FF0EF;
mem['h02EB] = 32'h1B448593;
mem['h02EC] = 32'h00040513;
mem['h02ED] = 32'hDBCFF0EF;
mem['h02EE] = 32'h00000693;
mem['h02EF] = 32'h00400593;
mem['h02F0] = 32'h00DA0633;
mem['h02F1] = 32'h026CC703;
mem['h02F2] = 32'h00064603;
mem['h02F3] = 32'h2CC70E63;
mem['h02F4] = 32'h40C70733;
mem['h02F5] = 32'h001AC683;
mem['h02F6] = 32'h26071263;
mem['h02F7] = 32'h02AAC603;
mem['h02F8] = 32'h00800713;
mem['h02F9] = 32'h24E61C63;
mem['h02FA] = 32'h02BAC703;
mem['h02FB] = 32'h24071863;
mem['h02FC] = 32'h004AAC83;
mem['h02FD] = 32'h00100713;
mem['h02FE] = 32'h00600613;
mem['h02FF] = 32'h80E18593;
mem['h0300] = 32'h610A8513;
mem['h0301] = 32'h60DA8423;
mem['h0302] = 32'h60EA85A3;
mem['h0303] = 32'h619AA623;
mem['h0304] = 32'hF38FF0EF;
mem['h0305] = 32'h00600613;
mem['h0306] = 32'h008A0593;
mem['h0307] = 32'h616A8513;
mem['h0308] = 32'hF28FF0EF;
mem['h0309] = 32'h00450737;
mem['h030A] = 32'h00870713;
mem['h030B] = 32'h60EAAE23;
mem['h030C] = 32'h018AD703;
mem['h030D] = 32'h00400613;
mem['h030E] = 32'h00090593;
mem['h030F] = 32'h62EA9023;
mem['h0310] = 32'h62AA8513;
mem['h0311] = 32'h01FF0737;
mem['h0312] = 32'h62EAA223;
mem['h0313] = 32'h620A9123;
mem['h0314] = 32'h620A9423;
mem['h0315] = 32'hEF4FF0EF;
mem['h0316] = 32'h00400613;
mem['h0317] = 32'h022A8593;
mem['h0318] = 32'h62EA8513;
mem['h0319] = 32'hEE4FF0EF;
mem['h031A] = 32'h01400593;
mem['h031B] = 32'h61EA8513;
mem['h031C] = 32'hDBCFF0EF;
mem['h031D] = 32'h00851713;
mem['h031E] = 32'h00855513;
mem['h031F] = 32'h00A76733;
mem['h0320] = 32'h62EA9423;
mem['h0321] = 32'h02EAD703;
mem['h0322] = 32'hFD6C8613;
mem['h0323] = 32'h032A8593;
mem['h0324] = 32'h62EA9B23;
mem['h0325] = 32'h030AD703;
mem['h0326] = 32'h63AA8513;
mem['h0327] = 32'h620A9923;
mem['h0328] = 32'h62EA9C23;
mem['h0329] = 32'h620A9A23;
mem['h032A] = 32'hEA0FF0EF;
mem['h032B] = 32'h80E18793;
mem['h032C] = 32'h62478513;
mem['h032D] = 32'hFDEC8593;
mem['h032E] = 32'hD74FF0EF;
mem['h032F] = 32'h00C12583;
mem['h0330] = 32'h00851713;
mem['h0331] = 32'h00855513;
mem['h0332] = 32'h00A76733;
mem['h0333] = 32'h00040513;
mem['h0334] = 32'h62EA9A23;
mem['h0335] = 32'hE98FF0EF;
mem['h0336] = 32'h000015B7;
mem['h0337] = 32'h22458593;
mem['h0338] = 32'h00040513;
mem['h0339] = 32'hC8CFF0EF;
mem['h033A] = 32'h004AD583;
mem['h033B] = 32'h13C0006F;
mem['h033C] = 32'h000017B7;
mem['h033D] = 32'h1FC78593;
mem['h033E] = 32'h00040513;
mem['h033F] = 32'hC74FF0EF;
mem['h0340] = 32'h004AD583;
mem['h0341] = 32'h00040513;
mem['h0342] = 32'hB94FF0EF;
mem['h0343] = 32'h1B448593;
mem['h0344] = 32'h00040513;
mem['h0345] = 32'hC5CFF0EF;
mem['h0346] = 32'h017AC603;
mem['h0347] = 32'h00100693;
mem['h0348] = 32'h016AC703;
mem['h0349] = 32'h10D61C63;
mem['h034A] = 32'h018AC683;
mem['h034B] = 32'h11A69863;
mem['h034C] = 32'h019AC683;
mem['h034D] = 32'h00D76733;
mem['h034E] = 32'h10071263;
mem['h034F] = 32'h00000693;
mem['h0350] = 32'h00400593;
mem['h0351] = 32'h00DA0633;
mem['h0352] = 32'h02ECC703;
mem['h0353] = 32'h00064603;
mem['h0354] = 32'h14C70263;
mem['h0355] = 32'h40C70733;
mem['h0356] = 32'h001AC683;
mem['h0357] = 32'h0E071063;
mem['h0358] = 32'h01CAC703;
mem['h0359] = 32'h0C071C63;
mem['h035A] = 32'h01DAC703;
mem['h035B] = 32'h00100613;
mem['h035C] = 32'h0CC71663;
mem['h035D] = 32'h60EA85A3;
mem['h035E] = 32'h00600613;
mem['h035F] = 32'h02A00713;
mem['h0360] = 32'h81E18593;
mem['h0361] = 32'h610A8513;
mem['h0362] = 32'h60DA8423;
mem['h0363] = 32'h60EAA623;
mem['h0364] = 32'hDB8FF0EF;
mem['h0365] = 32'h008A0593;
mem['h0366] = 32'h00600613;
mem['h0367] = 32'h616A8513;
mem['h0368] = 32'hDA8FF0EF;
mem['h0369] = 32'h01000737;
mem['h036A] = 32'h60870713;
mem['h036B] = 32'h60EAAE23;
mem['h036C] = 32'h04060737;
mem['h036D] = 32'h100007B7;
mem['h036E] = 32'h00870713;
mem['h036F] = 32'h00878593;
mem['h0370] = 32'h62EAA023;
mem['h0371] = 32'h00600613;
mem['h0372] = 32'h20000713;
mem['h0373] = 32'h626A8513;
mem['h0374] = 32'h62EA9223;
mem['h0375] = 32'hD74FF0EF;
mem['h0376] = 32'h00400613;
mem['h0377] = 32'h00090593;
mem['h0378] = 32'h62CA8513;
mem['h0379] = 32'hD64FF0EF;
mem['h037A] = 32'h00600613;
mem['h037B] = 32'h81E18593;
mem['h037C] = 32'h630A8513;
mem['h037D] = 32'hD54FF0EF;
mem['h037E] = 32'h00400613;
mem['h037F] = 32'h024A8593;
mem['h0380] = 32'h636A8513;
mem['h0381] = 32'hD44FF0EF;
mem['h0382] = 32'h00812583;
mem['h0383] = 32'h00040513;
mem['h0384] = 32'hD5CFF0EF;
mem['h0385] = 32'h000015B7;
mem['h0386] = 32'h21058593;
mem['h0387] = 32'h00040513;
mem['h0388] = 32'hB50FF0EF;
mem['h0389] = 32'h60CAD583;
mem['h038A] = 32'h00040513;
mem['h038B] = 32'hA70FF0EF;
mem['h038C] = 32'h1B448593;
mem['h038D] = 32'h00040513;
mem['h038E] = 32'hB38FF0EF;
mem['h038F] = 32'h001AC683;
mem['h0390] = 32'h00100713;
mem['h0391] = 32'h06E69C63;
mem['h0392] = 32'h00200713;
mem['h0393] = 32'h00EA8023;
mem['h0394] = 32'h00DA81A3;
mem['h0395] = 32'h01898593;
mem['h0396] = 32'h00040513;
mem['h0397] = 32'hD10FF0EF;
mem['h0398] = 32'h00442703;
mem['h0399] = 32'h00072703;
mem['h039A] = 32'h00072703;
mem['h039B] = 32'h00072583;
mem['h039C] = 32'hB605D2E3;
mem['h039D] = 32'h0FF5F713;
mem['h039E] = 32'h01200693;
mem['h039F] = 32'hB4D70CE3;
mem['h03A0] = 32'h0FF5F593;
mem['h03A1] = 32'h00B10823;
mem['h03A2] = 32'h05659463;
mem['h03A3] = 32'h00010823;
mem['h03A4] = 32'hB45FF06F;
mem['h03A5] = 32'h00168693;
mem['h03A6] = 32'h001C8C93;
mem['h03A7] = 32'hEAB694E3;
mem['h03A8] = 32'h00000713;
mem['h03A9] = 32'hEB5FF06F;
mem['h03AA] = 32'h00168693;
mem['h03AB] = 32'h001C8C93;
mem['h03AC] = 32'hD0B698E3;
mem['h03AD] = 32'h00000713;
mem['h03AE] = 32'hD1DFF06F;
mem['h03AF] = 32'h00200613;
mem['h03B0] = 32'hFAC690E3;
mem['h03B1] = 32'h00EA8023;
mem['h03B2] = 32'h00EA81A3;
mem['h03B3] = 32'hF89FF06F;
mem['h03B4] = 32'h00000C93;
mem['h03B5] = 32'h01010C13;
mem['h03B6] = 32'h07758863;
mem['h03B7] = 32'h00800D13;
mem['h03B8] = 32'h07F00D93;
mem['h03B9] = 32'h01A58463;
mem['h03BA] = 32'h0FB59863;
mem['h03BB] = 32'h03905863;
mem['h03BC] = 32'h00800593;
mem['h03BD] = 32'h00040513;
mem['h03BE] = 32'h97CFF0EF;
mem['h03BF] = 32'h02000593;
mem['h03C0] = 32'h00040513;
mem['h03C1] = 32'h970FF0EF;
mem['h03C2] = 32'h00800593;
mem['h03C3] = 32'h00040513;
mem['h03C4] = 32'hFFFC0C13;
mem['h03C5] = 32'hFFFC8C93;
mem['h03C6] = 32'h95CFF0EF;
mem['h03C7] = 32'h00442603;
mem['h03C8] = 32'h00062603;
mem['h03C9] = 32'h00062603;
mem['h03CA] = 32'h00062583;
mem['h03CB] = 32'hFE05D8E3;
mem['h03CC] = 32'h01F00793;
mem['h03CD] = 32'h02FC8663;
mem['h03CE] = 32'h0FF5F593;
mem['h03CF] = 32'h00BC0023;
mem['h03D0] = 32'h03658063;
mem['h03D1] = 32'hFB7590E3;
mem['h03D2] = 32'h00D00593;
mem['h03D3] = 32'h00040513;
mem['h03D4] = 32'h924FF0EF;
mem['h03D5] = 32'h00A00593;
mem['h03D6] = 32'h00040513;
mem['h03D7] = 32'h918FF0EF;
mem['h03D8] = 32'h000C0023;
mem['h03D9] = 32'h0FFCFC93;
mem['h03DA] = 32'hA60C86E3;
mem['h03DB] = 32'h000015B7;
mem['h03DC] = 32'h00040513;
mem['h03DD] = 32'h23858593;
mem['h03DE] = 32'h9F8FF0EF;
mem['h03DF] = 32'h01010593;
mem['h03E0] = 32'h00040513;
mem['h03E1] = 32'h9ECFF0EF;
mem['h03E2] = 32'h1B448593;
mem['h03E3] = 32'h00040513;
mem['h03E4] = 32'h9E0FF0EF;
mem['h03E5] = 32'h000015B7;
mem['h03E6] = 32'h00040513;
mem['h03E7] = 32'h24458593;
mem['h03E8] = 32'h9D0FF0EF;
mem['h03E9] = 32'h000C8593;
mem['h03EA] = 32'h00040513;
mem['h03EB] = 32'h8F0FF0EF;
mem['h03EC] = 32'h1B448593;
mem['h03ED] = 32'h00040513;
mem['h03EE] = 32'h9B8FF0EF;
mem['h03EF] = 32'h01014583;
mem['h03F0] = 32'h00040513;
mem['h03F1] = 32'hB28FF0EF;
mem['h03F2] = 32'h1B448593;
mem['h03F3] = 32'h00040513;
mem['h03F4] = 32'h9A0FF0EF;
mem['h03F5] = 32'h9F9FF06F;
mem['h03F6] = 32'h00040513;
mem['h03F7] = 32'h898FF0EF;
mem['h03F8] = 32'h001C0C13;
mem['h03F9] = 32'h001C8C93;
mem['h03FA] = 32'hF35FF06F;
mem['h03FB] = 32'h06054063;
mem['h03FC] = 32'h0605C663;
mem['h03FD] = 32'h00058613;
mem['h03FE] = 32'h00050593;
mem['h03FF] = 32'hFFF00513;
mem['h0400] = 32'h02060C63;
mem['h0401] = 32'h00100693;
mem['h0402] = 32'h00B67A63;
mem['h0403] = 32'h00C05863;
mem['h0404] = 32'h00161613;
mem['h0405] = 32'h00169693;
mem['h0406] = 32'hFEB66AE3;
mem['h0407] = 32'h00000513;
mem['h0408] = 32'h00C5E663;
mem['h0409] = 32'h40C585B3;
mem['h040A] = 32'h00D56533;
mem['h040B] = 32'h0016D693;
mem['h040C] = 32'h00165613;
mem['h040D] = 32'hFE0696E3;
mem['h040E] = 32'h00008067;
mem['h040F] = 32'h00008293;
mem['h0410] = 32'hFB5FF0EF;
mem['h0411] = 32'h00058513;
mem['h0412] = 32'h00028067;
mem['h0413] = 32'h40A00533;
mem['h0414] = 32'h00B04863;
mem['h0415] = 32'h40B005B3;
mem['h0416] = 32'hF9DFF06F;
mem['h0417] = 32'h40B005B3;
mem['h0418] = 32'h00008293;
mem['h0419] = 32'hF91FF0EF;
mem['h041A] = 32'h40A00533;
mem['h041B] = 32'h00028067;
mem['h041C] = 32'h00008293;
mem['h041D] = 32'h0005CA63;
mem['h041E] = 32'h00054C63;
mem['h041F] = 32'hF79FF0EF;
mem['h0420] = 32'h00058513;
mem['h0421] = 32'h00028067;
mem['h0422] = 32'h40B005B3;
mem['h0423] = 32'hFE0558E3;
mem['h0424] = 32'h40A00533;
mem['h0425] = 32'hF61FF0EF;
mem['h0426] = 32'h40B00533;
mem['h0427] = 32'h00028067;
mem['h0428] = 32'h33323130;
mem['h0429] = 32'h37363534;
mem['h042A] = 32'h42413938;
mem['h042B] = 32'h46454443;
mem['h042C] = 32'h00000000;
mem['h042D] = 32'h3D3D3D3D;
mem['h042E] = 32'h3D3D3D3D;
mem['h042F] = 32'h3D3D3D3D;
mem['h0430] = 32'h3D3D3D3D;
mem['h0431] = 32'h3D3D3D3D;
mem['h0432] = 32'h3D3D3D3D;
mem['h0433] = 32'h3D3D3D3D;
mem['h0434] = 32'h3D3D3D3D;
mem['h0435] = 32'h3D3D3D3D;
mem['h0436] = 32'h3D3D3D3D;
mem['h0437] = 32'h0A0D3D3D;
mem['h0438] = 32'h00000000;
mem['h0439] = 32'h20202020;
mem['h043A] = 32'h57202020;
mem['h043B] = 32'h47657269;
mem['h043C] = 32'h64726175;
mem['h043D] = 32'h47504620;
mem['h043E] = 32'h79622041;
mem['h043F] = 32'h69684320;
mem['h0440] = 32'h6843696C;
mem['h0441] = 32'h20737069;
mem['h0442] = 32'h20202020;
mem['h0443] = 32'h0A0D2020;
mem['h0444] = 32'h00000000;
mem['h0445] = 32'h7774654E;
mem['h0446] = 32'h206B726F;
mem['h0447] = 32'h666E6F63;
mem['h0448] = 32'h72756769;
mem['h0449] = 32'h6F697461;
mem['h044A] = 32'h000A0D6E;
mem['h044B] = 32'h49202D2D;
mem['h044C] = 32'h64612050;
mem['h044D] = 32'h73657264;
mem['h044E] = 32'h20203A73;
mem['h044F] = 32'h20202020;
mem['h0450] = 32'h00002020;
mem['h0451] = 32'h2D2D0A0D;
mem['h0452] = 32'h62755320;
mem['h0453] = 32'h2074656E;
mem['h0454] = 32'h6B73616D;
mem['h0455] = 32'h2020203A;
mem['h0456] = 32'h20202020;
mem['h0457] = 32'h00000000;
mem['h0458] = 32'h2D2D0A0D;
mem['h0459] = 32'h43414D20;
mem['h045A] = 32'h64646120;
mem['h045B] = 32'h73736572;
mem['h045C] = 32'h2020203A;
mem['h045D] = 32'h20202020;
mem['h045E] = 32'h00000000;
mem['h045F] = 32'h2D2D0A0D;
mem['h0460] = 32'h66654420;
mem['h0461] = 32'h746C7561;
mem['h0462] = 32'h74616720;
mem['h0463] = 32'h79617765;
mem['h0464] = 32'h2020203A;
mem['h0465] = 32'h00000000;
mem['h0466] = 32'h2D2D0A0D;
mem['h0467] = 32'h66654420;
mem['h0468] = 32'h746C7561;
mem['h0469] = 32'h746E6920;
mem['h046A] = 32'h61667265;
mem['h046B] = 32'h203A6563;
mem['h046C] = 32'h00000000;
mem['h046D] = 32'h00000A0D;
mem['h046E] = 32'h2D2D2D2D;
mem['h046F] = 32'h2D2D2D2D;
mem['h0470] = 32'h2D2D2D2D;
mem['h0471] = 32'h2D2D2D2D;
mem['h0472] = 32'h2D2D2D2D;
mem['h0473] = 32'h2D2D2D2D;
mem['h0474] = 32'h2D2D2D2D;
mem['h0475] = 32'h2D2D2D2D;
mem['h0476] = 32'h2D2D2D2D;
mem['h0477] = 32'h2D2D2D2D;
mem['h0478] = 32'h0A0D2D2D;
mem['h0479] = 32'h00000000;
mem['h047A] = 32'h4E203C3C;
mem['h047B] = 32'h505F5445;
mem['h047C] = 32'h4F544F52;
mem['h047D] = 32'h4D43495F;
mem['h047E] = 32'h00203A50;
mem['h047F] = 32'h4E203C3C;
mem['h0480] = 32'h505F5445;
mem['h0481] = 32'h4F544F52;
mem['h0482] = 32'h5052415F;
mem['h0483] = 32'h0000203A;
mem['h0484] = 32'h4E203E3E;
mem['h0485] = 32'h505F5445;
mem['h0486] = 32'h4F544F52;
mem['h0487] = 32'h5052415F;
mem['h0488] = 32'h0000203A;
mem['h0489] = 32'h4E203E3E;
mem['h048A] = 32'h505F5445;
mem['h048B] = 32'h4F544F52;
mem['h048C] = 32'h4D43495F;
mem['h048D] = 32'h00203A50;
mem['h048E] = 32'h65636552;
mem['h048F] = 32'h64657669;
mem['h0490] = 32'h0000203A;
mem['h0491] = 32'h65636552;
mem['h0492] = 32'h64657669;
mem['h0493] = 32'h6E656C20;
mem['h0494] = 32'h3A687467;
mem['h0495] = 32'h00000020;
mem['h0496] = 32'h6301A8C0;
mem['h0497] = 32'h00FFFFFF;
mem['h0498] = 32'hAECCCACA;
mem['h0499] = 32'hA8C00100;
mem['h049A] = 32'h0001FE01;
mem['h049B] = 32'h00000000;
