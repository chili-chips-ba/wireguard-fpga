-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.9455399354105367]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 33
entity VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_1CLK_051b2cdc is
port(
 clk : in std_logic;
 elem_val : in unsigned(31 downto 0);
 ref_toks_0 : in chacha20_state;
 var_dim_0 : in unsigned(3 downto 0);
 return_output : out uint32_t_array_16_t);
end VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_1CLK_051b2cdc;
architecture arch of VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_1CLK_051b2cdc is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 1;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output : unsigned(31 downto 0);
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_return_output : unsigned(0 downto 0);

-- rv_data_15_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24]
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_cond : unsigned(0 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iftrue : unsigned(31 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iffalse : unsigned(31 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_return_output : unsigned(0 downto 0);

-- rv_data_12_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd]
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_cond : unsigned(0 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iftrue : unsigned(31 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iffalse : unsigned(31 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iftrue : unsigned(31 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iffalse : unsigned(31 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iftrue : unsigned(31 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iffalse : unsigned(31 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_return_output : unsigned(0 downto 0);

-- rv_data_10_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5]
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_cond : unsigned(0 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iftrue : unsigned(31 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iffalse : unsigned(31 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iftrue : unsigned(31 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iffalse : unsigned(31 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_return_output : unsigned(0 downto 0);

-- rv_data_13_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a]
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_cond : unsigned(0 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iftrue : unsigned(31 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iffalse : unsigned(31 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iftrue : unsigned(31 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iffalse : unsigned(31 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iftrue : unsigned(31 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iffalse : unsigned(31 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_return_output : unsigned(0 downto 0);

-- rv_data_8_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3]
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_cond : unsigned(0 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iftrue : unsigned(31 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iffalse : unsigned(31 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_return_output : unsigned(0 downto 0);

-- rv_data_11_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86]
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_cond : unsigned(0 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iftrue : unsigned(31 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iffalse : unsigned(31 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_return_output : unsigned(0 downto 0);

-- rv_data_14_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202]
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_cond : unsigned(0 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iftrue : unsigned(31 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iffalse : unsigned(31 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iftrue : unsigned(31 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iffalse : unsigned(31 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iftrue : unsigned(31 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iffalse : unsigned(31 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iftrue : unsigned(31 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iffalse : unsigned(31 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_return_output : unsigned(0 downto 0);

-- rv_data_9_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9]
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_cond : unsigned(0 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iftrue : unsigned(31 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iffalse : unsigned(31 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_return_output : unsigned(31 downto 0);

function CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_f407( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint32_t_array_16_t is
 
  variable base : uint32_t_array_16_t; 
  variable return_output : uint32_t_array_16_t;
begin
      base.data(15) := ref_toks_0;
      base.data(12) := ref_toks_1;
      base.data(1) := ref_toks_2;
      base.data(4) := ref_toks_3;
      base.data(10) := ref_toks_4;
      base.data(7) := ref_toks_5;
      base.data(13) := ref_toks_6;
      base.data(5) := ref_toks_7;
      base.data(2) := ref_toks_8;
      base.data(8) := ref_toks_9;
      base.data(11) := ref_toks_10;
      base.data(14) := ref_toks_11;
      base.data(3) := ref_toks_12;
      base.data(0) := ref_toks_13;
      base.data(6) := ref_toks_14;
      base.data(9) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_return_output);

-- rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24 : 1 clocks latency
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_cond,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iftrue,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iffalse,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_return_output);

-- rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd : 1 clocks latency
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_cond,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iftrue,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iffalse,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648 : 0 clocks latency
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934 : 1 clocks latency
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_return_output);

-- rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5 : 1 clocks latency
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_cond,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iftrue,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iffalse,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1 : 1 clocks latency
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_return_output);

-- rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a : 1 clocks latency
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_cond,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iftrue,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iffalse,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a : 1 clocks latency
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7 : 0 clocks latency
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_return_output);

-- rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3 : 1 clocks latency
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_cond,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iftrue,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iffalse,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_return_output);

-- rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86 : 1 clocks latency
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_cond,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iftrue,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iffalse,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_return_output);

-- rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202 : 1 clocks latency
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_cond,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iftrue,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iffalse,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560 : 0 clocks latency
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343 : 0 clocks latency
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7 : 1 clocks latency
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_return_output);

-- rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9 : 1 clocks latency
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_0b9cb19c port map (
clk,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_cond,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iftrue,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iffalse,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- Registers
 -- Stage 0
 REG_STAGE0_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output,
 REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output,
 REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output,
 REG_STAGE0_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_return_output,
 rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_return_output,
 rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_return_output,
 rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_return_output,
 rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_return_output,
 rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_return_output,
 rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_return_output,
 rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_return_output,
 rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(31 downto 0);
 variable VAR_ref_toks_0 : chacha20_state;
 variable VAR_var_dim_0 : unsigned(3 downto 0);
 variable VAR_return_output : uint32_t_array_16_t;
 variable VAR_base : chacha20_state;
 variable VAR_rv : uint32_t_array_16_t;
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c16_4097_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c16_1d7f_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c15_255d_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_d3a2_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_fd7a_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c15_c110_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c16_6d9d_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_7164_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_2afe_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c15_0f8d_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_03c8_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c16_5bad_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_3463_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c15_19f3_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c15_0241_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c15_d44f_return_output : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_f407_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_84d5_return_output : uint32_t_array_16_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_right := to_unsigned(14, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_right := to_unsigned(9, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_right := to_unsigned(12, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_right := to_unsigned(10, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_right := to_unsigned(8, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_right := to_unsigned(13, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_right := to_unsigned(11, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_right := to_unsigned(15, 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iftrue := VAR_elem_val;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iftrue := VAR_elem_val;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iftrue := VAR_elem_val;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iftrue := VAR_elem_val;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iftrue := VAR_elem_val;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iftrue := VAR_elem_val;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iftrue := VAR_elem_val;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iftrue := VAR_elem_val;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_left := VAR_var_dim_0;
     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c15_c110] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c15_c110_return_output := VAR_ref_toks_0.state(7);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_2afe] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_2afe_return_output := VAR_ref_toks_0.state(2);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_7164] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_7164_return_output := VAR_ref_toks_0.state(5);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c15_255d] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c15_255d_return_output := VAR_ref_toks_0.state(1);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c15_19f3] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c15_19f3_return_output := VAR_ref_toks_0.state(0);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c16_1d7f] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c16_1d7f_return_output := VAR_ref_toks_0.state(12);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c16_6d9d] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c16_6d9d_return_output := VAR_ref_toks_0.state(13);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_d3a2] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_d3a2_return_output := VAR_ref_toks_0.state(4);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c15_d44f] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c15_d44f_return_output := VAR_ref_toks_0.state(9);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_fd7a] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_fd7a_return_output := VAR_ref_toks_0.state(10);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c15_0f8d] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c15_0f8d_return_output := VAR_ref_toks_0.state(8);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c16_5bad] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c16_5bad_return_output := VAR_ref_toks_0.state(14);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_03c8] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_03c8_return_output := VAR_ref_toks_0.state(11);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c16_4097] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c16_4097_return_output := VAR_ref_toks_0.state(15);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_3463] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_3463_return_output := VAR_ref_toks_0.state(3);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c15_0241] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c15_0241_return_output := VAR_ref_toks_0.state(6);

     -- Submodule level 1
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_3d46_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_4ea6_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_51e6_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_2418_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_e291_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_835b_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_aa70_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_a6f1_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_2db4_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_53cc_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_c1b9_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_4092_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_b38a_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_f4b8_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_6d5b_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7b0e_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c15_19f3_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_fd7a_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_03c8_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c16_1d7f_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c16_6d9d_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c16_5bad_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c16_4097_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c15_255d_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_2afe_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_3463_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_d3a2_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_7164_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c15_0241_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c15_c110_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c15_0f8d_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c15_d44f_return_output;
     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a] LATENCY=1
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_iffalse;

     -- rv_data_9_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9] LATENCY=1
     -- Inputs
     rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_cond <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_cond;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iftrue <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iftrue;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iffalse <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_iffalse;

     -- rv_data_8_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3] LATENCY=1
     -- Inputs
     rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_cond <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_cond;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iftrue <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iftrue;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iffalse <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_iffalse;

     -- rv_data_11_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86] LATENCY=1
     -- Inputs
     rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_cond <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_cond;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iftrue <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iftrue;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iffalse <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_iffalse;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934] LATENCY=1
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_iffalse;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1] LATENCY=1
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_iffalse;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7] LATENCY=1
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_iffalse;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output;

     -- rv_data_12_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd] LATENCY=1
     -- Inputs
     rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_cond <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_cond;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iftrue <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iftrue;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iffalse <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_iffalse;

     -- rv_data_14_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202] LATENCY=1
     -- Inputs
     rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_cond <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_cond;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iftrue <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iftrue;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iffalse <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_iffalse;

     -- rv_data_13_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a] LATENCY=1
     -- Inputs
     rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_cond <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_cond;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iftrue <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iftrue;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iffalse <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_iffalse;

     -- rv_data_15_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24] LATENCY=1
     -- Inputs
     rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_cond <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_cond;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iftrue <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iftrue;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iffalse <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_iffalse;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output;

     -- rv_data_10_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5] LATENCY=1
     -- Inputs
     rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_cond <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_cond;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iftrue <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iftrue;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iffalse <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_iffalse;

     -- Submodule level 2
     -- Write to comb signals
     COMB_STAGE0_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output;
     COMB_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output;
     COMB_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output;
     COMB_STAGE0_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output := REG_STAGE0_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output := REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output := REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output := REG_STAGE0_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output;
     -- Submodule outputs
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_return_output := rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_return_output := rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_return_output := rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_return_output := rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_return_output := rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_return_output := rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_return_output := rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_return_output := rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_return_output;

     -- Submodule level 0
     -- CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_f407[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_84d5] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_f407_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_84d5_return_output := CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_f407(
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_bb24_return_output,
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_43cd_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_4934_return_output,
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_37f5_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_d5c1_return_output,
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_733a_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_732a_return_output,
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output,
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_83d3_return_output,
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_0d86_return_output,
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_7202_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_d0d7_return_output,
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_a8c9_return_output);

     -- Submodule level 1
     VAR_return_output := VAR_CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_f407_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_84d5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     REG_STAGE0_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output <= COMB_STAGE0_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_2648_return_output;
     REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output <= COMB_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_7ba7_return_output;
     REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output <= COMB_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_3560_return_output;
     REG_STAGE0_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output <= COMB_STAGE0_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_1343_return_output;
 end if;
end process;

end arch;
