-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 16
entity axis128_keep_count_0CLK_08de2a73 is
port(
 axis : in axis128_t;
 return_output : out unsigned(4 downto 0));
end axis128_keep_count_0CLK_08de2a73;
architecture arch of axis128_keep_count_0CLK_08de2a73 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS[axis_h_l91_c5_4225]
signal FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS[axis_h_l91_c5_ce9a]
signal FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS[axis_h_l91_c5_ffe3]
signal FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS[axis_h_l91_c5_a61e]
signal FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS[axis_h_l91_c5_f944]
signal FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS[axis_h_l91_c5_942b]
signal FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS[axis_h_l91_c5_65be]
signal FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS[axis_h_l91_c5_536d]
signal FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS[axis_h_l91_c5_d52c]
signal FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS[axis_h_l91_c5_a7a8]
signal FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS[axis_h_l91_c5_1a72]
signal FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS[axis_h_l91_c5_df26]
signal FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS[axis_h_l91_c5_86a4]
signal FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS[axis_h_l91_c5_667e]
signal FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS[axis_h_l91_c5_81f1]
signal FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS[axis_h_l91_c5_5012]
signal FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_return_output : unsigned(5 downto 0);


begin

-- SUBMODULE INSTANCES 
-- FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225 : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_left,
FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_right,
FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_left,
FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_right,
FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3 : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_left,
FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_right,
FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_left,
FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_right,
FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944 : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_left,
FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_right,
FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_left,
FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_right,
FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_left,
FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_right,
FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_left,
FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_right,
FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_left,
FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_right,
FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8 : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_left,
FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_right,
FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72 : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_left,
FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_right,
FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26 : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_left,
FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_right,
FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4 : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_left,
FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_right,
FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_left,
FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_right,
FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1 : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_left,
FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_right,
FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_return_output);

-- FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012 : 0 clocks latency
FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_left,
FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_right,
FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 axis,
 -- All submodule outputs
 FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_return_output,
 FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(4 downto 0);
 variable VAR_axis : axis128_t;
 variable VAR_rv : unsigned(4 downto 0);
 variable VAR_i : unsigned(31 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_rv_axis_h_l91_c5_5fc4 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_bf29_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_return_output : unsigned(5 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_left := to_unsigned(0, 5);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_axis := axis;

     -- Submodule level 0
     -- FOR_axis_h_l90_c3_f6b2_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(11);

     -- FOR_axis_h_l90_c3_f6b2_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(0);

     -- FOR_axis_h_l90_c3_f6b2_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(15);

     -- FOR_axis_h_l90_c3_f6b2_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(10);

     -- FOR_axis_h_l90_c3_f6b2_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(4);

     -- FOR_axis_h_l90_c3_f6b2_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(14);

     -- FOR_axis_h_l90_c3_f6b2_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(5);

     -- FOR_axis_h_l90_c3_f6b2_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(8);

     -- FOR_axis_h_l90_c3_f6b2_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(3);

     -- FOR_axis_h_l90_c3_f6b2_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(13);

     -- FOR_axis_h_l90_c3_f6b2_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(9);

     -- FOR_axis_h_l90_c3_f6b2_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(12);

     -- FOR_axis_h_l90_c3_f6b2_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(2);

     -- FOR_axis_h_l90_c3_f6b2_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(7);

     -- FOR_axis_h_l90_c3_f6b2_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(6);

     -- FOR_axis_h_l90_c3_f6b2_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d[axis_h_l91_c11_bf29] LATENCY=0
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_bf29_return_output := VAR_axis.tkeep(1);

     -- Submodule level 1
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_bf29_return_output;
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_right := VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_bf29_return_output;
     -- FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS[axis_h_l91_c5_4225] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_left;
     FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_return_output := FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_return_output;

     -- Submodule level 2
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_4225_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_0_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS[axis_h_l91_c5_ce9a] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_left;
     FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_return_output := FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_return_output;

     -- Submodule level 3
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ce9a_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_1_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS[axis_h_l91_c5_ffe3] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_left;
     FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_return_output := FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_return_output;

     -- Submodule level 4
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_ffe3_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_2_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS[axis_h_l91_c5_a61e] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_left;
     FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_return_output := FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_return_output;

     -- Submodule level 5
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_a61e_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_3_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS[axis_h_l91_c5_f944] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_left;
     FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_return_output := FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_return_output;

     -- Submodule level 6
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_f944_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_4_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS[axis_h_l91_c5_942b] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_left;
     FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_return_output := FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_return_output;

     -- Submodule level 7
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_942b_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_5_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS[axis_h_l91_c5_65be] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_left;
     FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_return_output := FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_return_output;

     -- Submodule level 8
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_65be_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_6_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS[axis_h_l91_c5_536d] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_left;
     FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_return_output := FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_return_output;

     -- Submodule level 9
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_536d_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_7_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS[axis_h_l91_c5_d52c] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_left;
     FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_return_output := FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_return_output;

     -- Submodule level 10
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_d52c_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_8_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS[axis_h_l91_c5_a7a8] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_left;
     FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_return_output := FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_return_output;

     -- Submodule level 11
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_a7a8_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_9_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS[axis_h_l91_c5_1a72] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_left;
     FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_return_output := FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_return_output;

     -- Submodule level 12
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_1a72_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_10_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS[axis_h_l91_c5_df26] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_left;
     FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_return_output := FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_return_output;

     -- Submodule level 13
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_df26_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_11_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS[axis_h_l91_c5_86a4] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_left;
     FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_return_output := FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_return_output;

     -- Submodule level 14
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_86a4_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_12_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS[axis_h_l91_c5_667e] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_left;
     FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_return_output := FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_return_output;

     -- Submodule level 15
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_667e_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_13_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS[axis_h_l91_c5_81f1] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_left;
     FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_return_output := FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_return_output;

     -- Submodule level 16
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_81f1_return_output, 5);
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_left := VAR_FOR_axis_h_l90_c3_f6b2_ITER_14_rv_axis_h_l91_c5_5fc4;
     -- FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS[axis_h_l91_c5_5012] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_left <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_left;
     FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_right <= VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_return_output := FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_return_output;

     -- Submodule level 17
     VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_rv_axis_h_l91_c5_5fc4 := resize(VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_5012_return_output, 5);
     VAR_return_output := VAR_FOR_axis_h_l90_c3_f6b2_ITER_15_rv_axis_h_l91_c5_5fc4;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
