-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 27
entity chacha20_block_0CLK_f1a496f6 is
port(
 state : in chacha20_state;
 return_output : out chacha20_state);
end chacha20_block_0CLK_f1a496f6;
architecture arch of chacha20_block_0CLK_f1a496f6 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- chacha20_block_step[chacha20_h_l72_c28_fcf3]
signal chacha20_block_step_chacha20_h_l72_c28_fcf3_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l72_c28_fcf3_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l73_c28_378a]
signal chacha20_block_step_chacha20_h_l73_c28_378a_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l73_c28_378a_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l74_c28_f57e]
signal chacha20_block_step_chacha20_h_l74_c28_f57e_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l74_c28_f57e_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l75_c28_e58f]
signal chacha20_block_step_chacha20_h_l75_c28_e58f_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l75_c28_e58f_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l76_c28_4b87]
signal chacha20_block_step_chacha20_h_l76_c28_4b87_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l76_c28_4b87_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l77_c28_1296]
signal chacha20_block_step_chacha20_h_l77_c28_1296_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l77_c28_1296_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l78_c28_ff0e]
signal chacha20_block_step_chacha20_h_l78_c28_ff0e_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l78_c28_ff0e_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l79_c28_873d]
signal chacha20_block_step_chacha20_h_l79_c28_873d_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l79_c28_873d_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l80_c28_2731]
signal chacha20_block_step_chacha20_h_l80_c28_2731_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l80_c28_2731_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l81_c29_1e3c]
signal chacha20_block_step_chacha20_h_l81_c29_1e3c_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output : chacha20_state;

-- FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS[chacha20_h_l87_c27_8a29]
signal FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);

function CONST_REF_RD_chacha20_state_chacha20_state_23da( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return chacha20_state is
 
  variable base : chacha20_state; 
  variable return_output : chacha20_state;
begin
      base.state(0) := ref_toks_0;
      base.state(1) := ref_toks_1;
      base.state(2) := ref_toks_2;
      base.state(3) := ref_toks_3;
      base.state(4) := ref_toks_4;
      base.state(5) := ref_toks_5;
      base.state(6) := ref_toks_6;
      base.state(7) := ref_toks_7;
      base.state(8) := ref_toks_8;
      base.state(9) := ref_toks_9;
      base.state(10) := ref_toks_10;
      base.state(11) := ref_toks_11;
      base.state(12) := ref_toks_12;
      base.state(13) := ref_toks_13;
      base.state(14) := ref_toks_14;
      base.state(15) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- chacha20_block_step_chacha20_h_l72_c28_fcf3 : 0 clocks latency
chacha20_block_step_chacha20_h_l72_c28_fcf3 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l72_c28_fcf3_state0,
chacha20_block_step_chacha20_h_l72_c28_fcf3_return_output);

-- chacha20_block_step_chacha20_h_l73_c28_378a : 0 clocks latency
chacha20_block_step_chacha20_h_l73_c28_378a : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l73_c28_378a_state0,
chacha20_block_step_chacha20_h_l73_c28_378a_return_output);

-- chacha20_block_step_chacha20_h_l74_c28_f57e : 0 clocks latency
chacha20_block_step_chacha20_h_l74_c28_f57e : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l74_c28_f57e_state0,
chacha20_block_step_chacha20_h_l74_c28_f57e_return_output);

-- chacha20_block_step_chacha20_h_l75_c28_e58f : 0 clocks latency
chacha20_block_step_chacha20_h_l75_c28_e58f : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l75_c28_e58f_state0,
chacha20_block_step_chacha20_h_l75_c28_e58f_return_output);

-- chacha20_block_step_chacha20_h_l76_c28_4b87 : 0 clocks latency
chacha20_block_step_chacha20_h_l76_c28_4b87 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l76_c28_4b87_state0,
chacha20_block_step_chacha20_h_l76_c28_4b87_return_output);

-- chacha20_block_step_chacha20_h_l77_c28_1296 : 0 clocks latency
chacha20_block_step_chacha20_h_l77_c28_1296 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l77_c28_1296_state0,
chacha20_block_step_chacha20_h_l77_c28_1296_return_output);

-- chacha20_block_step_chacha20_h_l78_c28_ff0e : 0 clocks latency
chacha20_block_step_chacha20_h_l78_c28_ff0e : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l78_c28_ff0e_state0,
chacha20_block_step_chacha20_h_l78_c28_ff0e_return_output);

-- chacha20_block_step_chacha20_h_l79_c28_873d : 0 clocks latency
chacha20_block_step_chacha20_h_l79_c28_873d : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l79_c28_873d_state0,
chacha20_block_step_chacha20_h_l79_c28_873d_return_output);

-- chacha20_block_step_chacha20_h_l80_c28_2731 : 0 clocks latency
chacha20_block_step_chacha20_h_l80_c28_2731 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l80_c28_2731_state0,
chacha20_block_step_chacha20_h_l80_c28_2731_return_output);

-- chacha20_block_step_chacha20_h_l81_c29_1e3c : 0 clocks latency
chacha20_block_step_chacha20_h_l81_c29_1e3c : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l81_c29_1e3c_state0,
chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);

-- FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : 0 clocks latency
FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29 : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left,
FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right,
FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 state,
 -- All submodule outputs
 chacha20_block_step_chacha20_h_l72_c28_fcf3_return_output,
 chacha20_block_step_chacha20_h_l73_c28_378a_return_output,
 chacha20_block_step_chacha20_h_l74_c28_f57e_return_output,
 chacha20_block_step_chacha20_h_l75_c28_e58f_return_output,
 chacha20_block_step_chacha20_h_l76_c28_4b87_return_output,
 chacha20_block_step_chacha20_h_l77_c28_1296_return_output,
 chacha20_block_step_chacha20_h_l78_c28_ff0e_return_output,
 chacha20_block_step_chacha20_h_l79_c28_873d_return_output,
 chacha20_block_step_chacha20_h_l80_c28_2731_return_output,
 chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output,
 FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : chacha20_state;
 variable VAR_state : chacha20_state;
 variable VAR_output : chacha20_state;
 variable VAR_step1 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l72_c28_fcf3_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l72_c28_fcf3_return_output : chacha20_state;
 variable VAR_step2 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l73_c28_378a_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l73_c28_378a_return_output : chacha20_state;
 variable VAR_step3 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l74_c28_f57e_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l74_c28_f57e_return_output : chacha20_state;
 variable VAR_step4 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l75_c28_e58f_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l75_c28_e58f_return_output : chacha20_state;
 variable VAR_step5 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l76_c28_4b87_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l76_c28_4b87_return_output : chacha20_state;
 variable VAR_step6 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l77_c28_1296_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l77_c28_1296_return_output : chacha20_state;
 variable VAR_step7 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l78_c28_ff0e_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l78_c28_ff0e_return_output : chacha20_state;
 variable VAR_step8 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l79_c28_873d_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l79_c28_873d_return_output : chacha20_state;
 variable VAR_step9 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l80_c28_2731_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l80_c28_2731_return_output : chacha20_state;
 variable VAR_step10 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output : chacha20_state;
 variable VAR_i : unsigned(3 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_output_state_0_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_output_state_1_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_output_state_2_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_output_state_3_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_output_state_4_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_output_state_5_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_output_state_6_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_output_state_7_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_output_state_8_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_output_state_9_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_output_state_10_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_output_state_11_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_output_state_12_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_output_state_13_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_output_state_14_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_output_state_15_chacha20_h_l87_c9_9f67 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c27_c979_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c45_f670_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output : unsigned(32 downto 0);
 variable VAR_CONST_REF_RD_chacha20_state_chacha20_state_23da_chacha20_h_l90_c12_6a92_return_output : chacha20_state;
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_state := state;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l72_c28_fcf3_state0 := VAR_state;
     -- FOR_chacha20_h_l85_c5_d0eb_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(7);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(2);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(9);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(4);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(3);

     -- chacha20_block_step[chacha20_h_l72_c28_fcf3] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l72_c28_fcf3_state0 <= VAR_chacha20_block_step_chacha20_h_l72_c28_fcf3_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l72_c28_fcf3_return_output := chacha20_block_step_chacha20_h_l72_c28_fcf3_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(11);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(14);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(5);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(6);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(1);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(8);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(10);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(15);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(13);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(0);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[chacha20_h_l87_c45_f670] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c45_f670_return_output := VAR_state.state(12);

     -- Submodule level 1
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c45_f670_return_output;
     VAR_chacha20_block_step_chacha20_h_l73_c28_378a_state0 := VAR_chacha20_block_step_chacha20_h_l72_c28_fcf3_return_output;
     -- chacha20_block_step[chacha20_h_l73_c28_378a] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l73_c28_378a_state0 <= VAR_chacha20_block_step_chacha20_h_l73_c28_378a_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l73_c28_378a_return_output := chacha20_block_step_chacha20_h_l73_c28_378a_return_output;

     -- Submodule level 2
     VAR_chacha20_block_step_chacha20_h_l74_c28_f57e_state0 := VAR_chacha20_block_step_chacha20_h_l73_c28_378a_return_output;
     -- chacha20_block_step[chacha20_h_l74_c28_f57e] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l74_c28_f57e_state0 <= VAR_chacha20_block_step_chacha20_h_l74_c28_f57e_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l74_c28_f57e_return_output := chacha20_block_step_chacha20_h_l74_c28_f57e_return_output;

     -- Submodule level 3
     VAR_chacha20_block_step_chacha20_h_l75_c28_e58f_state0 := VAR_chacha20_block_step_chacha20_h_l74_c28_f57e_return_output;
     -- chacha20_block_step[chacha20_h_l75_c28_e58f] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l75_c28_e58f_state0 <= VAR_chacha20_block_step_chacha20_h_l75_c28_e58f_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l75_c28_e58f_return_output := chacha20_block_step_chacha20_h_l75_c28_e58f_return_output;

     -- Submodule level 4
     VAR_chacha20_block_step_chacha20_h_l76_c28_4b87_state0 := VAR_chacha20_block_step_chacha20_h_l75_c28_e58f_return_output;
     -- chacha20_block_step[chacha20_h_l76_c28_4b87] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l76_c28_4b87_state0 <= VAR_chacha20_block_step_chacha20_h_l76_c28_4b87_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l76_c28_4b87_return_output := chacha20_block_step_chacha20_h_l76_c28_4b87_return_output;

     -- Submodule level 5
     VAR_chacha20_block_step_chacha20_h_l77_c28_1296_state0 := VAR_chacha20_block_step_chacha20_h_l76_c28_4b87_return_output;
     -- chacha20_block_step[chacha20_h_l77_c28_1296] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l77_c28_1296_state0 <= VAR_chacha20_block_step_chacha20_h_l77_c28_1296_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l77_c28_1296_return_output := chacha20_block_step_chacha20_h_l77_c28_1296_return_output;

     -- Submodule level 6
     VAR_chacha20_block_step_chacha20_h_l78_c28_ff0e_state0 := VAR_chacha20_block_step_chacha20_h_l77_c28_1296_return_output;
     -- chacha20_block_step[chacha20_h_l78_c28_ff0e] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l78_c28_ff0e_state0 <= VAR_chacha20_block_step_chacha20_h_l78_c28_ff0e_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l78_c28_ff0e_return_output := chacha20_block_step_chacha20_h_l78_c28_ff0e_return_output;

     -- Submodule level 7
     VAR_chacha20_block_step_chacha20_h_l79_c28_873d_state0 := VAR_chacha20_block_step_chacha20_h_l78_c28_ff0e_return_output;
     -- chacha20_block_step[chacha20_h_l79_c28_873d] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l79_c28_873d_state0 <= VAR_chacha20_block_step_chacha20_h_l79_c28_873d_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l79_c28_873d_return_output := chacha20_block_step_chacha20_h_l79_c28_873d_return_output;

     -- Submodule level 8
     VAR_chacha20_block_step_chacha20_h_l80_c28_2731_state0 := VAR_chacha20_block_step_chacha20_h_l79_c28_873d_return_output;
     -- chacha20_block_step[chacha20_h_l80_c28_2731] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l80_c28_2731_state0 <= VAR_chacha20_block_step_chacha20_h_l80_c28_2731_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l80_c28_2731_return_output := chacha20_block_step_chacha20_h_l80_c28_2731_return_output;

     -- Submodule level 9
     VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_state0 := VAR_chacha20_block_step_chacha20_h_l80_c28_2731_return_output;
     -- chacha20_block_step[chacha20_h_l81_c29_1e3c] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l81_c29_1e3c_state0 <= VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output := chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output;

     -- Submodule level 10
     -- FOR_chacha20_h_l85_c5_d0eb_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(11);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(7);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(4);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(3);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(2);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(1);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(14);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(15);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(12);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(9);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(8);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(10);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(6);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(13);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(5);

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[chacha20_h_l87_c27_c979] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c27_c979_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_1e3c_return_output.state(0);

     -- Submodule level 11
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c27_c979_return_output;
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left := VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c27_c979_return_output;
     -- FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS[chacha20_h_l87_c27_8a29] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_left;
     FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right <= VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output := FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output;

     -- Submodule level 12
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_output_state_0_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_output_state_10_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_output_state_11_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_output_state_12_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_output_state_13_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_output_state_14_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_output_state_15_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_output_state_1_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_output_state_2_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_output_state_3_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_output_state_4_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_output_state_5_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_output_state_6_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_output_state_7_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_output_state_8_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_output_state_9_chacha20_h_l87_c9_9f67 := resize(VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_8a29_return_output, 32);
     -- CONST_REF_RD_chacha20_state_chacha20_state_23da[chacha20_h_l90_c12_6a92] LATENCY=0
     VAR_CONST_REF_RD_chacha20_state_chacha20_state_23da_chacha20_h_l90_c12_6a92_return_output := CONST_REF_RD_chacha20_state_chacha20_state_23da(
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_0_output_state_0_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_1_output_state_1_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_2_output_state_2_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_3_output_state_3_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_4_output_state_4_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_5_output_state_5_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_6_output_state_6_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_7_output_state_7_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_8_output_state_8_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_9_output_state_9_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_10_output_state_10_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_11_output_state_11_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_12_output_state_12_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_13_output_state_13_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_14_output_state_14_chacha20_h_l87_c9_9f67,
     VAR_FOR_chacha20_h_l85_c5_d0eb_ITER_15_output_state_15_chacha20_h_l87_c9_9f67);

     -- Submodule level 13
     VAR_return_output := VAR_CONST_REF_RD_chacha20_state_chacha20_state_23da_chacha20_h_l90_c12_6a92_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
