mem['h0000] = 32'h00000093;
mem['h0001] = 32'h00000193;
mem['h0002] = 32'h00000213;
mem['h0003] = 32'h00000293;
mem['h0004] = 32'h00000313;
mem['h0005] = 32'h00000393;
mem['h0006] = 32'h00000413;
mem['h0007] = 32'h00000493;
mem['h0008] = 32'h00000513;
mem['h0009] = 32'h00000593;
mem['h000A] = 32'h00000613;
mem['h000B] = 32'h00000693;
mem['h000C] = 32'h00000713;
mem['h000D] = 32'h00000793;
mem['h000E] = 32'h00000813;
mem['h000F] = 32'h00000893;
mem['h0010] = 32'h00000913;
mem['h0011] = 32'h00000993;
mem['h0012] = 32'h00000A13;
mem['h0013] = 32'h00000A93;
mem['h0014] = 32'h00000B13;
mem['h0015] = 32'h00000B93;
mem['h0016] = 32'h00000C13;
mem['h0017] = 32'h00000C93;
mem['h0018] = 32'h00000D13;
mem['h0019] = 32'h00000D93;
mem['h001A] = 32'h00000E13;
mem['h001B] = 32'h00000E93;
mem['h001C] = 32'h00000F13;
mem['h001D] = 32'h00000F93;
mem['h001E] = 32'h00000517;
mem['h001F] = 32'h13050513;
mem['h0020] = 32'h00000593;
mem['h0021] = 32'h00000613;
mem['h0022] = 32'h00C5DC63;
mem['h0023] = 32'h00052683;
mem['h0024] = 32'h00D5A023;
mem['h0025] = 32'h00450513;
mem['h0026] = 32'h00458593;
mem['h0027] = 32'hFEC5C8E3;
mem['h0028] = 32'h00000513;
mem['h0029] = 32'h00000593;
mem['h002A] = 32'h00B55863;
mem['h002B] = 32'h00052023;
mem['h002C] = 32'h00450513;
mem['h002D] = 32'hFEB54CE3;
mem['h002E] = 32'h04C000EF;
mem['h002F] = 32'h0000006F;
mem['h0030] = 32'hFD010113;
mem['h0031] = 32'h02812623;
mem['h0032] = 32'h03010413;
mem['h0033] = 32'hFCA42E23;
mem['h0034] = 32'hFE042623;
mem['h0035] = 32'h0100006F;
mem['h0036] = 32'hFEC42783;
mem['h0037] = 32'h00178793;
mem['h0038] = 32'hFEF42623;
mem['h0039] = 32'hFEC42783;
mem['h003A] = 32'hFDC42703;
mem['h003B] = 32'hFEE7E6E3;
mem['h003C] = 32'h00000013;
mem['h003D] = 32'h00000013;
mem['h003E] = 32'h02C12403;
mem['h003F] = 32'h03010113;
mem['h0040] = 32'h00008067;
mem['h0041] = 32'hFE010113;
mem['h0042] = 32'h00112E23;
mem['h0043] = 32'h00812C23;
mem['h0044] = 32'h02010413;
mem['h0045] = 32'h200007B7;
mem['h0046] = 32'hFEF42623;
mem['h0047] = 32'hFEC42783;
mem['h0048] = 32'h0517C703;
mem['h0049] = 32'h00276713;
mem['h004A] = 32'h04E788A3;
mem['h004B] = 32'hFEC42783;
mem['h004C] = 32'h0507C783;
mem['h004D] = 32'h0017F793;
mem['h004E] = 32'h0FF7F713;
mem['h004F] = 32'hFEC42783;
mem['h0050] = 32'h00177713;
mem['h0051] = 32'h0517C683;
mem['h0052] = 32'hFFE6F693;
mem['h0053] = 32'h00E6E733;
mem['h0054] = 32'h04E788A3;
mem['h0055] = 32'h000F47B7;
mem['h0056] = 32'h24078513;
mem['h0057] = 32'hF65FF0EF;
mem['h0058] = 32'hFEC42783;
mem['h0059] = 32'h0517C703;
mem['h005A] = 32'hFFD77713;
mem['h005B] = 32'h04E788A3;
mem['h005C] = 32'hFEC42783;
mem['h005D] = 32'h0507C783;
mem['h005E] = 32'h0017F793;
mem['h005F] = 32'h0FF7F713;
mem['h0060] = 32'hFEC42783;
mem['h0061] = 32'h00177713;
mem['h0062] = 32'h0517C683;
mem['h0063] = 32'hFFE6F693;
mem['h0064] = 32'h00E6E733;
mem['h0065] = 32'h04E788A3;
mem['h0066] = 32'h000F47B7;
mem['h0067] = 32'h24078513;
mem['h0068] = 32'hF21FF0EF;
mem['h0069] = 32'hF79FF06F;
