-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 96
entity uint320_mul_0CLK_babc4282 is
port(
 a : in u320_t;
 b : in u320_t;
 return_output : out u320_t);
end uint320_mul_0CLK_babc4282;
architecture arch of uint320_mul_0CLK_babc4282 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_f673]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_888b]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_7942]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_0060]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_3a51]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_a228]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_6223]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_f05b]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_4823]
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_726a]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_d20d]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_e119]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_aee7]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_de62]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_9ae6]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_5198]
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_becb]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_dcb1]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_69ae]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_cb24]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_8d97]
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_92a7]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l132_c21_de68]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_a24b]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_6887]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l134_c22_7e98]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_11d9]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_bd9e]
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd]
signal FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2]
signal FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_6eb7]
signal FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_return_output : unsigned(64 downto 0);

function CONST_REF_RD_u320_t_u320_t_4216( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned) return u320_t is
 
  variable base : u320_t; 
  variable return_output : u320_t;
begin
      base.limbs(0) := ref_toks_0;
      base.limbs(1) := ref_toks_1;
      base.limbs(2) := ref_toks_2;
      base.limbs(3) := ref_toks_3;
      base.limbs(4) := ref_toks_4;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_left,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_right,
FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_left,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_right,
FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_left,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_right,
FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_left,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_right,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_left,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_right,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_left,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_right,
FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left,
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right,
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left,
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right,
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output);

-- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7 : 0 clocks latency
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_left,
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_right,
FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 a,
 b,
 -- All submodule outputs
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output,
 FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : u320_t;
 variable VAR_a : u320_t;
 variable VAR_b : u320_t;
 variable VAR_temp : u320_t;
 variable VAR_i : signed(31 downto 0);
 variable VAR_carry : unsigned(63 downto 0);
 variable VAR_j : signed(31 downto 0);
 variable VAR_high : unsigned(63 downto 0);
 variable VAR_low : unsigned(63 downto 0);
 variable VAR_product : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_old_value : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_8c38_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_8c38_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_8c38_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_8c38_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_d752_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_8c38_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_8121_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_return_output : unsigned(64 downto 0);
 variable VAR_res : u320_t;
 variable VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_5f71_return_output : u320_t;
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_8121_DUPLICATE_8da0_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_d752_DUPLICATE_146f_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_d752_DUPLICATE_3d28_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_d752_DUPLICATE_bd21_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_d752_DUPLICATE_6274_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_8121_DUPLICATE_4834_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_8121_DUPLICATE_bfd1_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_8121_DUPLICATE_f7e0_return_output : unsigned(63 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue := to_unsigned(1, 1);
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l128_c34_8c38] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_8c38_return_output := u320_t_NULL.limbs(4);

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l128_c34_8c38] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_8c38_return_output := u320_t_NULL.limbs(3);

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l128_c34_8c38] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_8c38_return_output := u320_t_NULL.limbs(1);

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l128_c34_8c38] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_8c38_return_output := u320_t_NULL.limbs(0);

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l128_c34_8c38] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_8c38_return_output := u320_t_NULL.limbs(2);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_8c38_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_8c38_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_8c38_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_8c38_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_8c38_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_a := a;
     VAR_b := b;

     -- Submodule level 0
     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c32_8121]_DUPLICATE_f7e0 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_8121_DUPLICATE_f7e0_return_output := VAR_a.limbs(3);

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c45_d752] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_d752_return_output := VAR_b.limbs(4);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c32_8121]_DUPLICATE_bfd1 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_8121_DUPLICATE_bfd1_return_output := VAR_a.limbs(2);

     -- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c32_8121] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_8121_return_output := VAR_a.limbs(4);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c45_d752]_DUPLICATE_146f LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_d752_DUPLICATE_146f_return_output := VAR_b.limbs(0);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c45_d752]_DUPLICATE_3d28 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_d752_DUPLICATE_3d28_return_output := VAR_b.limbs(1);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c45_d752]_DUPLICATE_bd21 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_d752_DUPLICATE_bd21_return_output := VAR_b.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c45_d752]_DUPLICATE_6274 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_d752_DUPLICATE_6274_return_output := VAR_b.limbs(3);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c32_8121]_DUPLICATE_8da0 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_8121_DUPLICATE_8da0_return_output := VAR_a.limbs(0);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c32_8121]_DUPLICATE_4834 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_8121_DUPLICATE_4834_return_output := VAR_a.limbs(1);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_8121_DUPLICATE_8da0_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_8121_DUPLICATE_8da0_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_8121_DUPLICATE_8da0_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_8121_DUPLICATE_8da0_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_8121_DUPLICATE_8da0_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_d752_DUPLICATE_146f_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_d752_DUPLICATE_146f_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_d752_DUPLICATE_146f_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_d752_DUPLICATE_146f_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_d752_DUPLICATE_146f_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_8121_DUPLICATE_4834_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_8121_DUPLICATE_4834_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_8121_DUPLICATE_4834_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_8121_DUPLICATE_4834_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_d752_DUPLICATE_3d28_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_d752_DUPLICATE_3d28_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_d752_DUPLICATE_3d28_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_d752_DUPLICATE_3d28_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_8121_DUPLICATE_bfd1_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_8121_DUPLICATE_bfd1_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_8121_DUPLICATE_bfd1_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_d752_DUPLICATE_bd21_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_d752_DUPLICATE_bd21_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_d752_DUPLICATE_bd21_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_8121_DUPLICATE_f7e0_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_8121_DUPLICATE_f7e0_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_d752_DUPLICATE_6274_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_d752_DUPLICATE_6274_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_d752_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_8121_return_output;
     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_09bd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_09bd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_product_poly1305_h_l127_c22_282d_0;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_product_poly1305_h_l127_c22_282d_0;
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_f673] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- Submodule level 4
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f673_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output;

     -- Submodule level 5
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l132_c21_de68_return_output;
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- Submodule level 6
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output;
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_888b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_return_output;

     -- Submodule level 7
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_888b_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a;
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_7942] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_return_output;

     -- Submodule level 8
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_7942_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- Submodule level 9
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_726a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_return_output;

     -- Submodule level 10
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_726a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_0060] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_return_output;

     -- Submodule level 11
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0060_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a;
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_3a51] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- Submodule level 12
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3a51_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_d20d] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_return_output;

     -- Submodule level 13
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d20d_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_e119] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_return_output;

     -- Submodule level 14
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e119_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_a228] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- Submodule level 15
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a228_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_2_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_becb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_6223] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_return_output;

     -- Submodule level 16
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_6223_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_becb_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l133_c13_1176;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l133_c13_1176;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_aee7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_return_output;

     -- Submodule level 17
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_aee7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_de62] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- Submodule level 18
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_MUX_poly1305_h_l134_c22_7e98_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de62_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_f05b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_dcb1] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- Submodule level 19
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_f05b_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l132_c21_de68_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_dcb1_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_3_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_4823] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_left;
     FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_return_output := FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_69ae] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_return_output;

     -- Submodule level 20
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4823_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_MUX_poly1305_h_l134_c22_7e98_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_69ae_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_4_low_poly1305_h_l133_c13_1176;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_9ae6] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output;

     -- Submodule level 21
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_9ae6_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l132_c21_de68_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_2_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_a24b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_left;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_92a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_5198] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_left;
     FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_return_output := FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- Submodule level 22
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_5198_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_MUX_poly1305_h_l134_c22_7e98_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_92a7_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_a24b_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_3_low_poly1305_h_l133_c13_1176;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l132_c21_de68] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_cb24] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_6887] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_left;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;

     -- Submodule level 23
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_cb24_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_6887_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l132_c21_de68_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_1_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX[poly1305_h_l134_c22_7e98] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_cond;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iftrue;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_8d97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_left;
     FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_return_output := FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_return_output;

     -- Submodule level 24
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8d97_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_MUX_poly1305_h_l134_c22_7e98_return_output;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_2_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_11d9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_left;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_return_output;

     -- Submodule level 25
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_11d9_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_high_poly1305_h_l134_c13_2e2a;
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_bd9e] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_left;
     FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_return_output := FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_return_output;

     -- Submodule level 26
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_bd9e_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right := VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_1_low_poly1305_h_l133_c13_1176;
     -- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_f1c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_left;
     FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output := FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output;

     -- Submodule level 27
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_f1c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_left := VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l131_c13_b045;
     -- FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_6eb7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_left <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_left;
     FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_right <= VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_return_output := FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_return_output;

     -- Submodule level 28
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176 := resize(VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6eb7_return_output, 64);
     -- CONST_REF_RD_u320_t_u320_t_4216[poly1305_h_l141_c18_5f71] LATENCY=0
     VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_5f71_return_output := CONST_REF_RD_u320_t_u320_t_4216(
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_0_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176,
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_1_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176,
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_2_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176,
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_3_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176,
     VAR_FOR_poly1305_h_l120_c5_0067_ITER_4_FOR_poly1305_h_l123_c9_6562_ITER_0_low_poly1305_h_l133_c13_1176);

     -- Submodule level 29
     VAR_return_output := VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_5f71_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
